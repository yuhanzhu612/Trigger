module InstFetch(
  input         clock,
  input         reset,
  output        io_imem_inst_valid,
  input         io_imem_inst_ready,
  output [31:0] io_imem_inst_addr,
  input  [31:0] io_imem_inst_read,
  output [31:0] io_fe_pc,
  output [31:0] io_fe_inst,
  input         io_br_valid,
  input         io_br_taken,
  input  [31:0] io_br_target,
  input         io_csr_jmp,
  input  [31:0] io_newpc,
  output        io_instr_valid,
  input         io_flush,
  output        io_if_valid_out,
  input         io_if_allow_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  if_valid_in; // @[InstFetch.scala 34:28]
  reg  abandon; // @[InstFetch.scala 39:30]
  reg  wait_valid; // @[InstFetch.scala 40:30]
  reg [31:0] wait_pc; // @[InstFetch.scala 41:30]
  wire  branch_valid = io_br_taken & io_br_valid; // @[InstFetch.scala 42:35]
  reg  flush_wait; // @[InstFetch.scala 44:27]
  reg  csr_jmp_wait; // @[InstFetch.scala 45:29]
  reg [31:0] csr_jmp_wait_pc; // @[InstFetch.scala 46:32]
  wire  csr_jmp = io_csr_jmp | csr_jmp_wait | flush_wait; // @[InstFetch.scala 47:44]
  wire [31:0] csr_newpc = io_csr_jmp ? io_newpc : csr_jmp_wait_pc; // @[InstFetch.scala 48:22]
  wire  hands_done = io_imem_inst_ready & io_imem_inst_valid; // @[InstFetch.scala 50:42]
  wire  _preif_ready_go_T_1 = ~wait_valid; // @[InstFetch.scala 52:51]
  wire  preif_ready_go = hands_done & ~wait_valid & ~csr_jmp_wait; // @[InstFetch.scala 52:63]
  wire  if_allow_in = ~if_valid_in | io_if_valid_out & io_if_allow_out; // @[InstFetch.scala 59:32]
  wire  _GEN_0 = if_allow_in ? preif_ready_go : if_valid_in; // @[InstFetch.scala 60:21 InstFetch.scala 61:17 InstFetch.scala 34:28]
  wire  _GEN_1 = io_imem_inst_ready ? 1'h0 : csr_jmp_wait; // @[InstFetch.scala 68:33 InstFetch.scala 69:18 InstFetch.scala 45:29]
  wire  _GEN_2 = io_csr_jmp | _GEN_1; // @[InstFetch.scala 64:21 InstFetch.scala 65:18]
  wire  _GEN_4 = io_imem_inst_ready ? 1'h0 : flush_wait; // @[InstFetch.scala 75:33 InstFetch.scala 76:16 InstFetch.scala 44:27]
  wire  _GEN_5 = csr_jmp_wait | _GEN_4; // @[InstFetch.scala 72:23 InstFetch.scala 73:16]
  wire  _GEN_6 = io_imem_inst_ready ? 1'h0 : wait_valid; // @[InstFetch.scala 83:33 InstFetch.scala 84:16 InstFetch.scala 40:30]
  wire  _GEN_7 = branch_valid | _GEN_6; // @[InstFetch.scala 79:23 InstFetch.scala 80:16]
  wire  _GEN_9 = io_imem_inst_ready ? 1'h0 : abandon; // @[InstFetch.scala 90:33 InstFetch.scala 91:13 InstFetch.scala 39:30]
  wire  _GEN_10 = wait_valid | _GEN_9; // @[InstFetch.scala 87:21 InstFetch.scala 88:13]
  reg [31:0] if_pc; // @[InstFetch.scala 94:22]
  reg [31:0] if_inst; // @[InstFetch.scala 95:24]
  wire [31:0] _next_pc_T_2 = if_pc + 32'h4; // @[InstFetch.scala 96:115]
  wire [31:0] _next_pc_T_3 = wait_valid | abandon ? wait_pc : _next_pc_T_2; // @[InstFetch.scala 96:76]
  wire [31:0] _next_pc_T_4 = branch_valid ? io_br_target : _next_pc_T_3; // @[InstFetch.scala 96:44]
  assign io_imem_inst_valid = ~if_valid_in | io_if_valid_out & io_if_allow_out; // @[InstFetch.scala 59:32]
  assign io_imem_inst_addr = csr_jmp ? csr_newpc : _next_pc_T_4; // @[InstFetch.scala 96:20]
  assign io_fe_pc = io_flush ? 32'h0 : if_pc; // @[InstFetch.scala 119:21]
  assign io_fe_inst = io_flush ? 32'h0 : if_inst; // @[InstFetch.scala 120:21]
  assign io_instr_valid = io_flush ? 1'h0 : 1'h1; // @[InstFetch.scala 126:24]
  assign io_if_valid_out = if_valid_in & _preif_ready_go_T_1; // @[InstFetch.scala 57:31]
  always @(posedge clock) begin
    if_valid_in <= reset | _GEN_0; // @[InstFetch.scala 34:28 InstFetch.scala 34:28]
    if (reset) begin // @[InstFetch.scala 39:30]
      abandon <= 1'h0; // @[InstFetch.scala 39:30]
    end else begin
      abandon <= _GEN_10;
    end
    if (reset) begin // @[InstFetch.scala 40:30]
      wait_valid <= 1'h0; // @[InstFetch.scala 40:30]
    end else begin
      wait_valid <= _GEN_7;
    end
    if (reset) begin // @[InstFetch.scala 41:30]
      wait_pc <= 32'h0; // @[InstFetch.scala 41:30]
    end else if (branch_valid) begin // @[InstFetch.scala 79:23]
      wait_pc <= io_br_target; // @[InstFetch.scala 81:13]
    end
    if (reset) begin // @[InstFetch.scala 44:27]
      flush_wait <= 1'h0; // @[InstFetch.scala 44:27]
    end else begin
      flush_wait <= _GEN_5;
    end
    if (reset) begin // @[InstFetch.scala 45:29]
      csr_jmp_wait <= 1'h0; // @[InstFetch.scala 45:29]
    end else begin
      csr_jmp_wait <= _GEN_2;
    end
    if (reset) begin // @[InstFetch.scala 46:32]
      csr_jmp_wait_pc <= 32'h0; // @[InstFetch.scala 46:32]
    end else if (io_csr_jmp) begin // @[InstFetch.scala 48:22]
      csr_jmp_wait_pc <= io_newpc;
    end
    if (reset) begin // @[InstFetch.scala 94:22]
      if_pc <= 32'h7ffffffc; // @[InstFetch.scala 94:22]
    end else if (if_allow_in & preif_ready_go) begin // @[InstFetch.scala 109:41]
      if (io_flush) begin // @[InstFetch.scala 110:19]
        if_pc <= 32'h0;
      end else if (csr_jmp) begin // @[InstFetch.scala 96:20]
        if_pc <= csr_newpc;
      end else begin
        if_pc <= _next_pc_T_4;
      end
    end
    if (reset) begin // @[InstFetch.scala 95:24]
      if_inst <= 32'h0; // @[InstFetch.scala 95:24]
    end else if (if_allow_in & preif_ready_go) begin // @[InstFetch.scala 109:41]
      if (io_flush) begin // @[InstFetch.scala 111:19]
        if_inst <= 32'h0;
      end else begin
        if_inst <= io_imem_inst_read;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  if_valid_in = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  abandon = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wait_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  wait_pc = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  flush_wait = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  csr_jmp_wait = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  csr_jmp_wait_pc = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  if_pc = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  if_inst = _RAND_8[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decode(
  input         clock,
  input         reset,
  output [4:0]  io_rs1_addr,
  output        io_rs1_en,
  input  [63:0] io_rs1_data,
  output [4:0]  io_rs2_addr,
  output        io_rs2_en,
  input  [63:0] io_rs2_data,
  input  [31:0] io_fe_pc,
  input  [31:0] io_fe_inst,
  output [31:0] io_id_pc,
  output [31:0] io_id_inst,
  output        io_id_wen,
  output [4:0]  io_id_wdest,
  output [63:0] io_id_op1,
  output [63:0] io_id_op2,
  output [63:0] io_rs2_value,
  input         io_mem_stall,
  input         io_instr_valid,
  input         io_time_int,
  input  [4:0]  io_EX_wdest,
  input  [4:0]  io_WB_wdest,
  input  [63:0] io_EX_result,
  input  [63:0] io_WB_result,
  output        io_type_w,
  output [11:0] io_idop_aluop,
  output [6:0]  io_idop_loadop,
  output [3:0]  io_idop_storeop,
  output [3:0]  io_idop_sysop,
  output        io_inst_my,
  output        io_skip,
  output [63:0] io_print,
  output        io_br_valid,
  output        io_br_taken,
  output [31:0] io_br_target,
  output        io_br_stall,
  input         io_flush,
  output        io_if_allow_out,
  output        io_id_valid_out,
  input         io_if_valid_out,
  input         io_id_allow_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  id_valid_in; // @[Decode.scala 52:28]
  wire  id_allow_in = ~id_valid_in | io_id_valid_out & io_id_allow_out; // @[Decode.scala 62:29]
  reg [31:0] id_pc; // @[Decode.scala 65:25]
  reg [31:0] id_inst; // @[Decode.scala 66:25]
  reg  instr_valid; // @[Decode.scala 71:28]
  wire [51:0] imm_i_hi = id_inst[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [11:0] imm_i_lo = id_inst[31:20]; // @[Decode.scala 92:43]
  wire [63:0] imm_i = {imm_i_hi,imm_i_lo}; // @[Cat.scala 30:58]
  wire [31:0] imm_u_hi_hi = id_inst[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [19:0] imm_u_hi_lo = id_inst[31:12]; // @[Decode.scala 93:43]
  wire [63:0] imm_u = {imm_u_hi_hi,imm_u_hi_lo,12'h0}; // @[Cat.scala 30:58]
  wire [42:0] imm_j_hi_hi_hi = id_inst[31] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 72:12]
  wire [7:0] imm_j_hi_lo = id_inst[19:12]; // @[Decode.scala 94:53]
  wire  imm_j_lo_hi_hi = id_inst[20]; // @[Decode.scala 94:67]
  wire [9:0] imm_j_lo_hi_lo = id_inst[30:21]; // @[Decode.scala 94:77]
  wire [63:0] imm_j = {imm_j_hi_hi_hi,id_inst[31],imm_j_hi_lo,imm_j_lo_hi_hi,imm_j_lo_hi_lo,1'h0}; // @[Cat.scala 30:58]
  wire  imm_b_hi_lo = id_inst[7]; // @[Decode.scala 95:53]
  wire [5:0] imm_b_lo_hi_hi = id_inst[30:25]; // @[Decode.scala 95:62]
  wire [3:0] imm_b_lo_hi_lo = id_inst[11:8]; // @[Decode.scala 95:76]
  wire [55:0] imm_b = {imm_j_hi_hi_hi,id_inst[31],imm_b_hi_lo,imm_b_lo_hi_hi,imm_b_lo_hi_lo,1'h0}; // @[Cat.scala 30:58]
  wire [6:0] imm_s_hi_lo = id_inst[31:25]; // @[Decode.scala 96:43]
  wire [4:0] imm_s_lo = id_inst[11:7]; // @[Decode.scala 96:57]
  wire [63:0] imm_s = {imm_i_hi,imm_s_hi_lo,imm_s_lo}; // @[Cat.scala 30:58]
  wire  _rs1_forward_T = io_rs1_addr != 5'h0; // @[Decode.scala 111:34]
  wire  _rs1_forward_T_1 = io_rs1_addr == io_EX_wdest; // @[Decode.scala 111:59]
  wire  rs1_forward = io_rs1_addr != 5'h0 & (io_rs1_addr == io_EX_wdest | io_rs1_addr == io_WB_wdest) & io_rs1_en; // @[Decode.scala 111:107]
  wire  _rs2_forward_T = io_rs2_addr != 5'h0; // @[Decode.scala 112:34]
  wire  _rs2_forward_T_1 = io_rs2_addr == io_EX_wdest; // @[Decode.scala 112:59]
  wire  rs2_forward = io_rs2_addr != 5'h0 & (io_rs2_addr == io_EX_wdest | io_rs2_addr == io_WB_wdest) & io_rs2_en; // @[Decode.scala 112:107]
  wire [63:0] _rs1_value_T_1 = _rs1_forward_T_1 ? io_EX_result : io_WB_result; // @[Decode.scala 114:39]
  wire [63:0] rs1_value = rs1_forward ? _rs1_value_T_1 : io_rs1_data; // @[Decode.scala 114:22]
  wire [63:0] _rs2_value_T_1 = _rs2_forward_T_1 ? io_EX_result : io_WB_result; // @[Decode.scala 115:39]
  wire [63:0] rs2_value = rs2_forward ? _rs2_value_T_1 : io_rs2_data; // @[Decode.scala 115:22]
  wire [31:0] _T_1 = id_inst & 32'h707f; // @[Decode.scala 117:14]
  wire  _T_2 = 32'h13 == _T_1; // @[Decode.scala 117:14]
  wire [5:0] _GEN_6 = 32'h13 == _T_1 ? 6'h10 : 6'h0; // @[Decode.scala 117:24 Decode.scala 118:15]
  wire [11:0] _GEN_7 = 32'h13 == _T_1 ? 12'h1 : 12'h0; // @[Decode.scala 117:24 Decode.scala 119:15]
  wire [5:0] _GEN_10 = 32'h7013 == _T_1 ? 6'h10 : _GEN_6; // @[Decode.scala 125:24 Decode.scala 126:15]
  wire [11:0] _GEN_11 = 32'h7013 == _T_1 ? 12'h40 : _GEN_7; // @[Decode.scala 125:24 Decode.scala 127:15]
  wire  _GEN_12 = 32'h7013 == _T_1 | _T_2; // @[Decode.scala 125:24 Decode.scala 128:15]
  wire [5:0] _GEN_14 = 32'h4013 == _T_1 ? 6'h10 : _GEN_10; // @[Decode.scala 133:24 Decode.scala 134:15]
  wire [11:0] _GEN_15 = 32'h4013 == _T_1 ? 12'h10 : _GEN_11; // @[Decode.scala 133:24 Decode.scala 135:15]
  wire  _GEN_16 = 32'h4013 == _T_1 | _GEN_12; // @[Decode.scala 133:24 Decode.scala 136:15]
  wire [5:0] _GEN_18 = 32'h6013 == _T_1 ? 6'h10 : _GEN_14; // @[Decode.scala 141:23 Decode.scala 142:15]
  wire [11:0] _GEN_19 = 32'h6013 == _T_1 ? 12'h20 : _GEN_15; // @[Decode.scala 141:23 Decode.scala 143:15]
  wire  _GEN_20 = 32'h6013 == _T_1 | _GEN_16; // @[Decode.scala 141:23 Decode.scala 144:15]
  wire [31:0] _T_9 = id_inst & 32'hfc00707f; // @[Decode.scala 149:14]
  wire [5:0] _GEN_22 = 32'h1013 == _T_9 ? 6'h10 : _GEN_18; // @[Decode.scala 149:24 Decode.scala 150:15]
  wire [11:0] _GEN_23 = 32'h1013 == _T_9 ? 12'h80 : _GEN_19; // @[Decode.scala 149:24 Decode.scala 151:15]
  wire  _GEN_24 = 32'h1013 == _T_9 | _GEN_20; // @[Decode.scala 149:24 Decode.scala 152:15]
  wire [5:0] _GEN_26 = 32'h5013 == _T_9 ? 6'h10 : _GEN_22; // @[Decode.scala 157:24 Decode.scala 158:15]
  wire [11:0] _GEN_27 = 32'h5013 == _T_9 ? 12'h100 : _GEN_23; // @[Decode.scala 157:24 Decode.scala 159:15]
  wire  _GEN_28 = 32'h5013 == _T_9 | _GEN_24; // @[Decode.scala 157:24 Decode.scala 160:15]
  wire [5:0] _GEN_30 = 32'h40005013 == _T_9 ? 6'h10 : _GEN_26; // @[Decode.scala 165:24 Decode.scala 166:15]
  wire [11:0] _GEN_31 = 32'h40005013 == _T_9 ? 12'h200 : _GEN_27; // @[Decode.scala 165:24 Decode.scala 167:15]
  wire  _GEN_32 = 32'h40005013 == _T_9 | _GEN_28; // @[Decode.scala 165:24 Decode.scala 168:15]
  wire [5:0] _GEN_34 = 32'h2013 == _T_1 ? 6'h10 : _GEN_30; // @[Decode.scala 173:24 Decode.scala 174:15]
  wire [11:0] _GEN_35 = 32'h2013 == _T_1 ? 12'h4 : _GEN_31; // @[Decode.scala 173:24 Decode.scala 175:15]
  wire  _GEN_36 = 32'h2013 == _T_1 | _GEN_32; // @[Decode.scala 173:24 Decode.scala 176:15]
  wire [5:0] _GEN_38 = 32'h3013 == _T_1 ? 6'h10 : _GEN_34; // @[Decode.scala 181:25 Decode.scala 182:15]
  wire [11:0] _GEN_39 = 32'h3013 == _T_1 ? 12'h8 : _GEN_35; // @[Decode.scala 181:25 Decode.scala 183:15]
  wire  _GEN_40 = 32'h3013 == _T_1 | _GEN_36; // @[Decode.scala 181:25 Decode.scala 184:15]
  wire  _T_20 = 32'h1b == _T_1; // @[Decode.scala 189:14]
  wire [5:0] _GEN_42 = 32'h1b == _T_1 ? 6'h10 : _GEN_38; // @[Decode.scala 189:25 Decode.scala 190:15]
  wire [11:0] _GEN_43 = 32'h1b == _T_1 ? 12'h1 : _GEN_39; // @[Decode.scala 189:25 Decode.scala 191:15]
  wire  _GEN_44 = 32'h1b == _T_1 | _GEN_40; // @[Decode.scala 189:25 Decode.scala 192:15]
  wire [31:0] _T_21 = id_inst & 32'hfe00707f; // @[Decode.scala 198:14]
  wire [5:0] _GEN_47 = 32'h101b == _T_21 ? 6'h10 : _GEN_42; // @[Decode.scala 198:25 Decode.scala 199:15]
  wire [11:0] _GEN_48 = 32'h101b == _T_21 ? 12'h80 : _GEN_43; // @[Decode.scala 198:25 Decode.scala 200:15]
  wire  _GEN_49 = 32'h101b == _T_21 | _GEN_44; // @[Decode.scala 198:25 Decode.scala 201:15]
  wire  _GEN_51 = 32'h101b == _T_21 | _T_20; // @[Decode.scala 198:25 Decode.scala 204:15]
  wire [5:0] _GEN_52 = 32'h501b == _T_21 ? 6'h10 : _GEN_47; // @[Decode.scala 207:25 Decode.scala 208:15]
  wire [11:0] _GEN_53 = 32'h501b == _T_21 ? 12'h100 : _GEN_48; // @[Decode.scala 207:25 Decode.scala 209:15]
  wire  _GEN_54 = 32'h501b == _T_21 | _GEN_49; // @[Decode.scala 207:25 Decode.scala 210:15]
  wire  _GEN_56 = 32'h501b == _T_21 | _GEN_51; // @[Decode.scala 207:25 Decode.scala 213:15]
  wire [5:0] _GEN_57 = 32'h4000501b == _T_21 ? 6'h10 : _GEN_52; // @[Decode.scala 216:25 Decode.scala 217:15]
  wire [11:0] _GEN_58 = 32'h4000501b == _T_21 ? 12'h200 : _GEN_53; // @[Decode.scala 216:25 Decode.scala 218:15]
  wire  _GEN_59 = 32'h4000501b == _T_21 | _GEN_54; // @[Decode.scala 216:25 Decode.scala 219:15]
  wire  _GEN_61 = 32'h4000501b == _T_21 | _GEN_56; // @[Decode.scala 216:25 Decode.scala 222:15]
  wire  _T_28 = 32'h67 == _T_1; // @[Decode.scala 225:14]
  wire [63:0] _io_br_target_T_1 = rs1_value + imm_i; // @[Decode.scala 232:31]
  wire [5:0] _GEN_62 = 32'h67 == _T_1 ? 6'h2 : _GEN_57; // @[Decode.scala 225:24 Decode.scala 226:15]
  wire [11:0] _GEN_63 = 32'h67 == _T_1 ? 12'h1 : _GEN_58; // @[Decode.scala 225:24 Decode.scala 227:15]
  wire  _GEN_64 = 32'h67 == _T_1 | _GEN_59; // @[Decode.scala 225:24 Decode.scala 228:15]
  wire [63:0] _GEN_67 = 32'h67 == _T_1 ? _io_br_target_T_1 : 64'h0; // @[Decode.scala 225:24 Decode.scala 232:18 Decode.scala 109:16]
  wire [5:0] _GEN_68 = 32'h3 == _T_1 ? 6'h10 : _GEN_62; // @[Decode.scala 235:22 Decode.scala 236:15]
  wire [11:0] _GEN_69 = 32'h3 == _T_1 ? 12'h1 : _GEN_63; // @[Decode.scala 235:22 Decode.scala 237:15]
  wire  _GEN_70 = 32'h3 == _T_1 | _GEN_64; // @[Decode.scala 235:22 Decode.scala 238:15]
  wire [6:0] _GEN_72 = 32'h3 == _T_1 ? 7'h1 : 7'h0; // @[Decode.scala 235:22 Decode.scala 241:15]
  wire [5:0] _GEN_73 = 32'h4003 == _T_1 ? 6'h10 : _GEN_68; // @[Decode.scala 244:23 Decode.scala 245:15]
  wire [11:0] _GEN_74 = 32'h4003 == _T_1 ? 12'h1 : _GEN_69; // @[Decode.scala 244:23 Decode.scala 246:15]
  wire  _GEN_75 = 32'h4003 == _T_1 | _GEN_70; // @[Decode.scala 244:23 Decode.scala 247:15]
  wire [6:0] _GEN_77 = 32'h4003 == _T_1 ? 7'h2 : _GEN_72; // @[Decode.scala 244:23 Decode.scala 250:15]
  wire [5:0] _GEN_78 = 32'h1003 == _T_1 ? 6'h10 : _GEN_73; // @[Decode.scala 253:22 Decode.scala 254:15]
  wire [11:0] _GEN_79 = 32'h1003 == _T_1 ? 12'h1 : _GEN_74; // @[Decode.scala 253:22 Decode.scala 255:15]
  wire  _GEN_80 = 32'h1003 == _T_1 | _GEN_75; // @[Decode.scala 253:22 Decode.scala 256:15]
  wire [6:0] _GEN_82 = 32'h1003 == _T_1 ? 7'h4 : _GEN_77; // @[Decode.scala 253:22 Decode.scala 259:15]
  wire [5:0] _GEN_83 = 32'h5003 == _T_1 ? 6'h10 : _GEN_78; // @[Decode.scala 262:23 Decode.scala 263:15]
  wire [11:0] _GEN_84 = 32'h5003 == _T_1 ? 12'h1 : _GEN_79; // @[Decode.scala 262:23 Decode.scala 264:15]
  wire  _GEN_85 = 32'h5003 == _T_1 | _GEN_80; // @[Decode.scala 262:23 Decode.scala 265:15]
  wire [6:0] _GEN_87 = 32'h5003 == _T_1 ? 7'h8 : _GEN_82; // @[Decode.scala 262:23 Decode.scala 268:15]
  wire [5:0] _GEN_88 = 32'h2003 == _T_1 ? 6'h10 : _GEN_83; // @[Decode.scala 271:22 Decode.scala 272:15]
  wire [11:0] _GEN_89 = 32'h2003 == _T_1 ? 12'h1 : _GEN_84; // @[Decode.scala 271:22 Decode.scala 273:15]
  wire  _GEN_90 = 32'h2003 == _T_1 | _GEN_85; // @[Decode.scala 271:22 Decode.scala 274:15]
  wire [6:0] _GEN_92 = 32'h2003 == _T_1 ? 7'h10 : _GEN_87; // @[Decode.scala 271:22 Decode.scala 277:15]
  wire [5:0] _GEN_93 = 32'h6003 == _T_1 ? 6'h10 : _GEN_88; // @[Decode.scala 280:23 Decode.scala 281:15]
  wire [11:0] _GEN_94 = 32'h6003 == _T_1 ? 12'h1 : _GEN_89; // @[Decode.scala 280:23 Decode.scala 282:15]
  wire  _GEN_95 = 32'h6003 == _T_1 | _GEN_90; // @[Decode.scala 280:23 Decode.scala 283:15]
  wire [6:0] _GEN_97 = 32'h6003 == _T_1 ? 7'h20 : _GEN_92; // @[Decode.scala 280:23 Decode.scala 286:15]
  wire [5:0] _GEN_98 = 32'h3003 == _T_1 ? 6'h10 : _GEN_93; // @[Decode.scala 289:22 Decode.scala 290:15]
  wire [11:0] _GEN_99 = 32'h3003 == _T_1 ? 12'h1 : _GEN_94; // @[Decode.scala 289:22 Decode.scala 291:15]
  wire  _GEN_100 = 32'h3003 == _T_1 | _GEN_95; // @[Decode.scala 289:22 Decode.scala 292:15]
  wire [6:0] id_loadop = 32'h3003 == _T_1 ? 7'h40 : _GEN_97; // @[Decode.scala 289:22 Decode.scala 295:15]
  wire [5:0] _GEN_103 = 32'h2073 == _T_1 ? 6'h10 : _GEN_98; // @[Decode.scala 298:25 Decode.scala 299:15]
  wire [11:0] _GEN_104 = 32'h2073 == _T_1 ? 12'h1 : _GEN_99; // @[Decode.scala 298:25 Decode.scala 300:15]
  wire  _GEN_105 = 32'h2073 == _T_1 | _GEN_100; // @[Decode.scala 298:25 Decode.scala 301:15]
  wire [3:0] _GEN_107 = 32'h2073 == _T_1 ? 4'h2 : 4'h0; // @[Decode.scala 298:25 Decode.scala 304:14]
  wire [5:0] _GEN_108 = 32'h6073 == _T_1 ? 6'h10 : _GEN_103; // @[Decode.scala 307:26 Decode.scala 308:15]
  wire [11:0] _GEN_109 = 32'h6073 == _T_1 ? 12'h1 : _GEN_104; // @[Decode.scala 307:26 Decode.scala 309:15]
  wire  _GEN_110 = 32'h6073 == _T_1 | _GEN_105; // @[Decode.scala 307:26 Decode.scala 310:15]
  wire [3:0] _GEN_112 = 32'h6073 == _T_1 ? 4'h8 : _GEN_107; // @[Decode.scala 307:26 Decode.scala 313:14]
  wire [5:0] _GEN_113 = 32'h3073 == _T_1 ? 6'h10 : _GEN_108; // @[Decode.scala 316:25 Decode.scala 317:15]
  wire [11:0] _GEN_114 = 32'h3073 == _T_1 ? 12'h1 : _GEN_109; // @[Decode.scala 316:25 Decode.scala 318:15]
  wire  _GEN_115 = 32'h3073 == _T_1 | _GEN_110; // @[Decode.scala 316:25 Decode.scala 319:15]
  wire [3:0] _GEN_117 = 32'h3073 == _T_1 ? 4'h3 : _GEN_112; // @[Decode.scala 316:25 Decode.scala 322:14]
  wire [5:0] _GEN_118 = 32'h7073 == _T_1 ? 6'h10 : _GEN_113; // @[Decode.scala 325:26 Decode.scala 326:15]
  wire [11:0] _GEN_119 = 32'h7073 == _T_1 ? 12'h1 : _GEN_114; // @[Decode.scala 325:26 Decode.scala 327:15]
  wire  _GEN_120 = 32'h7073 == _T_1 | _GEN_115; // @[Decode.scala 325:26 Decode.scala 328:15]
  wire [3:0] _GEN_122 = 32'h7073 == _T_1 ? 4'h9 : _GEN_117; // @[Decode.scala 325:26 Decode.scala 331:14]
  wire [5:0] _GEN_123 = 32'h1073 == _T_1 ? 6'h10 : _GEN_118; // @[Decode.scala 334:25 Decode.scala 335:15]
  wire [11:0] _GEN_124 = 32'h1073 == _T_1 ? 12'h1 : _GEN_119; // @[Decode.scala 334:25 Decode.scala 336:15]
  wire  _GEN_125 = 32'h1073 == _T_1 | _GEN_120; // @[Decode.scala 334:25 Decode.scala 337:15]
  wire [3:0] _GEN_127 = 32'h1073 == _T_1 ? 4'h1 : _GEN_122; // @[Decode.scala 334:25 Decode.scala 340:14]
  wire [5:0] _GEN_128 = 32'h73 == id_inst ? 6'h10 : _GEN_123; // @[Decode.scala 343:25 Decode.scala 344:15]
  wire [11:0] _GEN_129 = 32'h73 == id_inst ? 12'h1 : _GEN_124; // @[Decode.scala 343:25 Decode.scala 345:15]
  wire  _GEN_130 = 32'h73 == id_inst ? 1'h0 : _GEN_125; // @[Decode.scala 343:25 Decode.scala 346:15]
  wire [3:0] _GEN_132 = 32'h73 == id_inst ? 4'h4 : _GEN_127; // @[Decode.scala 343:25 Decode.scala 349:14]
  wire  _T_56 = 32'h23 == _T_1; // @[Decode.scala 352:14]
  wire [5:0] _GEN_133 = 32'h23 == _T_1 ? 6'h4 : _GEN_128; // @[Decode.scala 352:22 Decode.scala 353:15]
  wire [11:0] _GEN_134 = 32'h23 == _T_1 ? 12'h1 : _GEN_129; // @[Decode.scala 352:22 Decode.scala 354:15]
  wire  _GEN_135 = 32'h23 == _T_1 | _GEN_130; // @[Decode.scala 352:22 Decode.scala 355:15]
  wire  _GEN_137 = 32'h23 == _T_1 ? 1'h0 : _GEN_130; // @[Decode.scala 352:22 Decode.scala 357:13]
  wire [3:0] _GEN_138 = 32'h23 == _T_1 ? 4'h1 : 4'h0; // @[Decode.scala 352:22 Decode.scala 358:16]
  wire [5:0] _GEN_139 = 32'h1023 == _T_1 ? 6'h4 : _GEN_133; // @[Decode.scala 361:22 Decode.scala 362:15]
  wire [11:0] _GEN_140 = 32'h1023 == _T_1 ? 12'h1 : _GEN_134; // @[Decode.scala 361:22 Decode.scala 363:15]
  wire  _GEN_141 = 32'h1023 == _T_1 | _GEN_135; // @[Decode.scala 361:22 Decode.scala 364:15]
  wire  _GEN_142 = 32'h1023 == _T_1 | _T_56; // @[Decode.scala 361:22 Decode.scala 365:15]
  wire  _GEN_143 = 32'h1023 == _T_1 ? 1'h0 : _GEN_137; // @[Decode.scala 361:22 Decode.scala 366:13]
  wire [3:0] _GEN_144 = 32'h1023 == _T_1 ? 4'h2 : _GEN_138; // @[Decode.scala 361:22 Decode.scala 367:16]
  wire [5:0] _GEN_145 = 32'h2023 == _T_1 ? 6'h4 : _GEN_139; // @[Decode.scala 370:22 Decode.scala 371:15]
  wire [11:0] _GEN_146 = 32'h2023 == _T_1 ? 12'h1 : _GEN_140; // @[Decode.scala 370:22 Decode.scala 372:15]
  wire  _GEN_147 = 32'h2023 == _T_1 | _GEN_141; // @[Decode.scala 370:22 Decode.scala 373:15]
  wire  _GEN_148 = 32'h2023 == _T_1 | _GEN_142; // @[Decode.scala 370:22 Decode.scala 374:15]
  wire  _GEN_149 = 32'h2023 == _T_1 ? 1'h0 : _GEN_143; // @[Decode.scala 370:22 Decode.scala 375:13]
  wire [3:0] _GEN_150 = 32'h2023 == _T_1 ? 4'h4 : _GEN_144; // @[Decode.scala 370:22 Decode.scala 376:16]
  wire [5:0] _GEN_151 = 32'h3023 == _T_1 ? 6'h4 : _GEN_145; // @[Decode.scala 379:22 Decode.scala 380:15]
  wire [11:0] _GEN_152 = 32'h3023 == _T_1 ? 12'h1 : _GEN_146; // @[Decode.scala 379:22 Decode.scala 381:15]
  wire  _GEN_153 = 32'h3023 == _T_1 | _GEN_147; // @[Decode.scala 379:22 Decode.scala 382:15]
  wire  _GEN_154 = 32'h3023 == _T_1 | _GEN_148; // @[Decode.scala 379:22 Decode.scala 383:15]
  wire  _GEN_155 = 32'h3023 == _T_1 ? 1'h0 : _GEN_149; // @[Decode.scala 379:22 Decode.scala 384:13]
  wire [3:0] id_storeop = 32'h3023 == _T_1 ? 4'h8 : _GEN_150; // @[Decode.scala 379:22 Decode.scala 385:16]
  wire [31:0] _T_63 = id_inst & 32'h7f; // @[Decode.scala 388:14]
  wire  _T_64 = 32'h17 == _T_63; // @[Decode.scala 388:14]
  wire [5:0] _GEN_157 = 32'h17 == _T_63 ? 6'h20 : _GEN_151; // @[Decode.scala 388:25 Decode.scala 389:15]
  wire [11:0] _GEN_158 = 32'h17 == _T_63 ? 12'h1 : _GEN_152; // @[Decode.scala 388:25 Decode.scala 390:15]
  wire  _GEN_159 = 32'h17 == _T_63 ? 1'h0 : _GEN_153; // @[Decode.scala 388:25 Decode.scala 391:15]
  wire  _GEN_160 = 32'h17 == _T_63 ? 1'h0 : _GEN_154; // @[Decode.scala 388:25 Decode.scala 392:15]
  wire  _GEN_161 = 32'h17 == _T_63 | _GEN_155; // @[Decode.scala 388:25 Decode.scala 393:15]
  wire [5:0] _GEN_162 = 32'h37 == _T_63 ? 6'h20 : _GEN_157; // @[Decode.scala 396:23 Decode.scala 397:15]
  wire [11:0] _GEN_163 = 32'h37 == _T_63 ? 12'h1 : _GEN_158; // @[Decode.scala 396:23 Decode.scala 398:15]
  wire  _GEN_164 = 32'h37 == _T_63 ? 1'h0 : _GEN_159; // @[Decode.scala 396:23 Decode.scala 399:15]
  wire  _GEN_165 = 32'h37 == _T_63 ? 1'h0 : _GEN_160; // @[Decode.scala 396:23 Decode.scala 400:15]
  wire  _GEN_166 = 32'h37 == _T_63 | _GEN_161; // @[Decode.scala 396:23 Decode.scala 401:15]
  wire [63:0] _GEN_304 = {{32'd0}, id_pc}; // @[Decode.scala 411:27]
  wire [63:0] _io_br_target_T_3 = _GEN_304 + imm_j; // @[Decode.scala 411:27]
  wire [5:0] _GEN_167 = 32'h6f == _T_63 ? 6'h2 : _GEN_162; // @[Decode.scala 404:23 Decode.scala 405:15]
  wire [11:0] _GEN_168 = 32'h6f == _T_63 ? 12'h1 : _GEN_163; // @[Decode.scala 404:23 Decode.scala 406:15]
  wire  _GEN_169 = 32'h6f == _T_63 ? 1'h0 : _GEN_164; // @[Decode.scala 404:23 Decode.scala 407:15]
  wire  _GEN_170 = 32'h6f == _T_63 ? 1'h0 : _GEN_165; // @[Decode.scala 404:23 Decode.scala 408:15]
  wire  _GEN_171 = 32'h6f == _T_63 | _GEN_166; // @[Decode.scala 404:23 Decode.scala 409:15]
  wire  _GEN_172 = 32'h6f == _T_63 | _T_28; // @[Decode.scala 404:23 Decode.scala 410:17]
  wire [63:0] _GEN_173 = 32'h6f == _T_63 ? _io_br_target_T_3 : _GEN_67; // @[Decode.scala 404:23 Decode.scala 411:18]
  wire [5:0] _GEN_174 = 32'h33 == _T_21 ? 6'h8 : _GEN_167; // @[Decode.scala 414:23 Decode.scala 415:15]
  wire [11:0] _GEN_175 = 32'h33 == _T_21 ? 12'h1 : _GEN_168; // @[Decode.scala 414:23 Decode.scala 416:15]
  wire  _GEN_176 = 32'h33 == _T_21 | _GEN_169; // @[Decode.scala 414:23 Decode.scala 417:15]
  wire  _GEN_177 = 32'h33 == _T_21 | _GEN_170; // @[Decode.scala 414:23 Decode.scala 418:15]
  wire  _GEN_178 = 32'h33 == _T_21 | _GEN_171; // @[Decode.scala 414:23 Decode.scala 419:15]
  wire [5:0] _GEN_179 = 32'h40000033 == _T_21 ? 6'h8 : _GEN_174; // @[Decode.scala 422:23 Decode.scala 423:15]
  wire [11:0] _GEN_180 = 32'h40000033 == _T_21 ? 12'h2 : _GEN_175; // @[Decode.scala 422:23 Decode.scala 424:15]
  wire  _GEN_181 = 32'h40000033 == _T_21 | _GEN_176; // @[Decode.scala 422:23 Decode.scala 425:15]
  wire  _GEN_182 = 32'h40000033 == _T_21 | _GEN_177; // @[Decode.scala 422:23 Decode.scala 426:15]
  wire  _GEN_183 = 32'h40000033 == _T_21 | _GEN_178; // @[Decode.scala 422:23 Decode.scala 427:15]
  wire [5:0] _GEN_184 = 32'h1033 == _T_21 ? 6'h8 : _GEN_179; // @[Decode.scala 430:23 Decode.scala 431:15]
  wire [11:0] _GEN_185 = 32'h1033 == _T_21 ? 12'h80 : _GEN_180; // @[Decode.scala 430:23 Decode.scala 432:15]
  wire  _GEN_186 = 32'h1033 == _T_21 | _GEN_181; // @[Decode.scala 430:23 Decode.scala 433:15]
  wire  _GEN_187 = 32'h1033 == _T_21 | _GEN_182; // @[Decode.scala 430:23 Decode.scala 434:15]
  wire  _GEN_188 = 32'h1033 == _T_21 | _GEN_183; // @[Decode.scala 430:23 Decode.scala 435:15]
  wire [5:0] _GEN_189 = 32'h2033 == _T_21 ? 6'h8 : _GEN_184; // @[Decode.scala 438:23 Decode.scala 439:15]
  wire [11:0] _GEN_190 = 32'h2033 == _T_21 ? 12'h4 : _GEN_185; // @[Decode.scala 438:23 Decode.scala 440:15]
  wire  _GEN_191 = 32'h2033 == _T_21 | _GEN_186; // @[Decode.scala 438:23 Decode.scala 441:15]
  wire  _GEN_192 = 32'h2033 == _T_21 | _GEN_187; // @[Decode.scala 438:23 Decode.scala 442:15]
  wire  _GEN_193 = 32'h2033 == _T_21 | _GEN_188; // @[Decode.scala 438:23 Decode.scala 443:15]
  wire [5:0] _GEN_194 = 32'h3033 == _T_21 ? 6'h8 : _GEN_189; // @[Decode.scala 446:24 Decode.scala 447:15]
  wire [11:0] _GEN_195 = 32'h3033 == _T_21 ? 12'h8 : _GEN_190; // @[Decode.scala 446:24 Decode.scala 448:15]
  wire  _GEN_196 = 32'h3033 == _T_21 | _GEN_191; // @[Decode.scala 446:24 Decode.scala 449:15]
  wire  _GEN_197 = 32'h3033 == _T_21 | _GEN_192; // @[Decode.scala 446:24 Decode.scala 450:15]
  wire  _GEN_198 = 32'h3033 == _T_21 | _GEN_193; // @[Decode.scala 446:24 Decode.scala 451:15]
  wire [5:0] _GEN_199 = 32'h4033 == _T_21 ? 6'h8 : _GEN_194; // @[Decode.scala 454:23 Decode.scala 455:15]
  wire [11:0] _GEN_200 = 32'h4033 == _T_21 ? 12'h10 : _GEN_195; // @[Decode.scala 454:23 Decode.scala 456:15]
  wire  _GEN_201 = 32'h4033 == _T_21 | _GEN_196; // @[Decode.scala 454:23 Decode.scala 457:15]
  wire  _GEN_202 = 32'h4033 == _T_21 | _GEN_197; // @[Decode.scala 454:23 Decode.scala 458:15]
  wire  _GEN_203 = 32'h4033 == _T_21 | _GEN_198; // @[Decode.scala 454:23 Decode.scala 459:15]
  wire [5:0] _GEN_204 = 32'h5033 == _T_21 ? 6'h8 : _GEN_199; // @[Decode.scala 462:23 Decode.scala 463:15]
  wire [11:0] _GEN_205 = 32'h5033 == _T_21 ? 12'h100 : _GEN_200; // @[Decode.scala 462:23 Decode.scala 464:15]
  wire  _GEN_206 = 32'h5033 == _T_21 | _GEN_201; // @[Decode.scala 462:23 Decode.scala 465:15]
  wire  _GEN_207 = 32'h5033 == _T_21 | _GEN_202; // @[Decode.scala 462:23 Decode.scala 466:15]
  wire  _GEN_208 = 32'h5033 == _T_21 | _GEN_203; // @[Decode.scala 462:23 Decode.scala 467:15]
  wire [5:0] _GEN_209 = 32'h40005033 == _T_21 ? 6'h8 : _GEN_204; // @[Decode.scala 470:23 Decode.scala 471:15]
  wire [11:0] _GEN_210 = 32'h40005033 == _T_21 ? 12'h200 : _GEN_205; // @[Decode.scala 470:23 Decode.scala 472:15]
  wire  _GEN_211 = 32'h40005033 == _T_21 | _GEN_206; // @[Decode.scala 470:23 Decode.scala 473:15]
  wire  _GEN_212 = 32'h40005033 == _T_21 | _GEN_207; // @[Decode.scala 470:23 Decode.scala 474:15]
  wire  _GEN_213 = 32'h40005033 == _T_21 | _GEN_208; // @[Decode.scala 470:23 Decode.scala 475:15]
  wire [5:0] _GEN_214 = 32'h6033 == _T_21 ? 6'h8 : _GEN_209; // @[Decode.scala 478:22 Decode.scala 479:15]
  wire [11:0] _GEN_215 = 32'h6033 == _T_21 ? 12'h20 : _GEN_210; // @[Decode.scala 478:22 Decode.scala 480:15]
  wire  _GEN_216 = 32'h6033 == _T_21 | _GEN_211; // @[Decode.scala 478:22 Decode.scala 481:15]
  wire  _GEN_217 = 32'h6033 == _T_21 | _GEN_212; // @[Decode.scala 478:22 Decode.scala 482:15]
  wire  _GEN_218 = 32'h6033 == _T_21 | _GEN_213; // @[Decode.scala 478:22 Decode.scala 483:15]
  wire [5:0] _GEN_219 = 32'h7033 == _T_21 ? 6'h8 : _GEN_214; // @[Decode.scala 486:23 Decode.scala 487:15]
  wire [11:0] _GEN_220 = 32'h7033 == _T_21 ? 12'h40 : _GEN_215; // @[Decode.scala 486:23 Decode.scala 488:15]
  wire  _GEN_221 = 32'h7033 == _T_21 | _GEN_216; // @[Decode.scala 486:23 Decode.scala 489:15]
  wire  _GEN_222 = 32'h7033 == _T_21 | _GEN_217; // @[Decode.scala 486:23 Decode.scala 490:15]
  wire  _GEN_223 = 32'h7033 == _T_21 | _GEN_218; // @[Decode.scala 486:23 Decode.scala 491:15]
  wire [5:0] _GEN_224 = 32'h3b == _T_21 ? 6'h8 : _GEN_219; // @[Decode.scala 494:24 Decode.scala 495:15]
  wire [11:0] _GEN_225 = 32'h3b == _T_21 ? 12'h1 : _GEN_220; // @[Decode.scala 494:24 Decode.scala 496:15]
  wire  _GEN_226 = 32'h3b == _T_21 | _GEN_221; // @[Decode.scala 494:24 Decode.scala 497:15]
  wire  _GEN_227 = 32'h3b == _T_21 | _GEN_222; // @[Decode.scala 494:24 Decode.scala 498:15]
  wire  _GEN_228 = 32'h3b == _T_21 | _GEN_223; // @[Decode.scala 494:24 Decode.scala 499:15]
  wire  _GEN_229 = 32'h3b == _T_21 | _GEN_61; // @[Decode.scala 494:24 Decode.scala 500:15]
  wire [5:0] _GEN_230 = 32'h4000003b == _T_21 ? 6'h8 : _GEN_224; // @[Decode.scala 503:24 Decode.scala 504:15]
  wire [11:0] _GEN_231 = 32'h4000003b == _T_21 ? 12'h2 : _GEN_225; // @[Decode.scala 503:24 Decode.scala 505:15]
  wire  _GEN_232 = 32'h4000003b == _T_21 | _GEN_226; // @[Decode.scala 503:24 Decode.scala 506:15]
  wire  _GEN_233 = 32'h4000003b == _T_21 | _GEN_227; // @[Decode.scala 503:24 Decode.scala 507:15]
  wire  _GEN_234 = 32'h4000003b == _T_21 | _GEN_228; // @[Decode.scala 503:24 Decode.scala 508:15]
  wire  _GEN_235 = 32'h4000003b == _T_21 | _GEN_229; // @[Decode.scala 503:24 Decode.scala 509:15]
  wire [5:0] _GEN_236 = 32'h103b == _T_21 ? 6'h8 : _GEN_230; // @[Decode.scala 512:24 Decode.scala 513:15]
  wire [11:0] _GEN_237 = 32'h103b == _T_21 ? 12'h80 : _GEN_231; // @[Decode.scala 512:24 Decode.scala 514:15]
  wire  _GEN_238 = 32'h103b == _T_21 | _GEN_232; // @[Decode.scala 512:24 Decode.scala 515:15]
  wire  _GEN_239 = 32'h103b == _T_21 | _GEN_233; // @[Decode.scala 512:24 Decode.scala 516:15]
  wire  _GEN_240 = 32'h103b == _T_21 | _GEN_234; // @[Decode.scala 512:24 Decode.scala 517:15]
  wire  _GEN_241 = 32'h103b == _T_21 | _GEN_235; // @[Decode.scala 512:24 Decode.scala 518:15]
  wire [5:0] _GEN_242 = 32'h503b == _T_21 ? 6'h8 : _GEN_236; // @[Decode.scala 521:24 Decode.scala 522:15]
  wire [11:0] _GEN_243 = 32'h503b == _T_21 ? 12'h100 : _GEN_237; // @[Decode.scala 521:24 Decode.scala 523:15]
  wire  _GEN_244 = 32'h503b == _T_21 | _GEN_238; // @[Decode.scala 521:24 Decode.scala 524:15]
  wire  _GEN_245 = 32'h503b == _T_21 | _GEN_239; // @[Decode.scala 521:24 Decode.scala 525:15]
  wire  _GEN_246 = 32'h503b == _T_21 | _GEN_240; // @[Decode.scala 521:24 Decode.scala 526:15]
  wire  _GEN_247 = 32'h503b == _T_21 | _GEN_241; // @[Decode.scala 521:24 Decode.scala 527:15]
  wire [5:0] _GEN_248 = 32'h4000503b == _T_21 ? 6'h8 : _GEN_242; // @[Decode.scala 530:24 Decode.scala 531:15]
  wire [11:0] _GEN_249 = 32'h4000503b == _T_21 ? 12'h200 : _GEN_243; // @[Decode.scala 530:24 Decode.scala 532:15]
  wire  _GEN_250 = 32'h4000503b == _T_21 | _GEN_244; // @[Decode.scala 530:24 Decode.scala 533:15]
  wire  _GEN_251 = 32'h4000503b == _T_21 | _GEN_245; // @[Decode.scala 530:24 Decode.scala 534:15]
  wire  _GEN_252 = 32'h4000503b == _T_21 | _GEN_246; // @[Decode.scala 530:24 Decode.scala 535:15]
  wire [5:0] _GEN_254 = 32'h30200073 == id_inst ? 6'h8 : _GEN_248; // @[Decode.scala 539:24 Decode.scala 540:15]
  wire [11:0] id_aluop = 32'h30200073 == id_inst ? 12'h200 : _GEN_249; // @[Decode.scala 539:24 Decode.scala 541:15]
  wire  _GEN_256 = 32'h30200073 == id_inst | _GEN_250; // @[Decode.scala 539:24 Decode.scala 542:15]
  wire  _GEN_257 = 32'h30200073 == id_inst | _GEN_251; // @[Decode.scala 539:24 Decode.scala 543:15]
  wire  _GEN_258 = 32'h30200073 == id_inst ? 1'h0 : _GEN_252; // @[Decode.scala 539:24 Decode.scala 544:15]
  wire [3:0] _GEN_259 = 32'h30200073 == id_inst ? 4'h5 : _GEN_132; // @[Decode.scala 539:24 Decode.scala 545:15]
  wire [63:0] _io_br_taken_T = rs1_forward ? _rs1_value_T_1 : io_rs1_data; // @[Decode.scala 553:40]
  wire [63:0] _io_br_taken_T_1 = rs2_forward ? _rs2_value_T_1 : io_rs2_data; // @[Decode.scala 553:63]
  wire [55:0] _GEN_305 = {{24'd0}, id_pc}; // @[Decode.scala 554:27]
  wire [55:0] _io_br_target_T_5 = _GEN_305 + imm_b; // @[Decode.scala 554:27]
  wire [5:0] _GEN_260 = 32'h63 == _T_1 ? 6'h1 : _GEN_254; // @[Decode.scala 548:23 Decode.scala 549:15]
  wire  _GEN_261 = 32'h63 == _T_1 | _GEN_256; // @[Decode.scala 548:23 Decode.scala 550:15]
  wire  _GEN_262 = 32'h63 == _T_1 | _GEN_257; // @[Decode.scala 548:23 Decode.scala 551:15]
  wire  _GEN_263 = 32'h63 == _T_1 ? 1'h0 : _GEN_258; // @[Decode.scala 548:23 Decode.scala 552:13]
  wire  _GEN_264 = 32'h63 == _T_1 ? $signed(_io_br_taken_T) == $signed(_io_br_taken_T_1) : _GEN_172; // @[Decode.scala 548:23 Decode.scala 553:17]
  wire [63:0] _GEN_265 = 32'h63 == _T_1 ? {{8'd0}, _io_br_target_T_5} : _GEN_173; // @[Decode.scala 548:23 Decode.scala 554:18]
  wire [5:0] _GEN_266 = 32'h1063 == _T_1 ? 6'h1 : _GEN_260; // @[Decode.scala 557:23 Decode.scala 558:15]
  wire  _GEN_267 = 32'h1063 == _T_1 | _GEN_261; // @[Decode.scala 557:23 Decode.scala 559:15]
  wire  _GEN_268 = 32'h1063 == _T_1 | _GEN_262; // @[Decode.scala 557:23 Decode.scala 560:15]
  wire  _GEN_269 = 32'h1063 == _T_1 ? 1'h0 : _GEN_263; // @[Decode.scala 557:23 Decode.scala 561:13]
  wire  _GEN_270 = 32'h1063 == _T_1 ? $signed(_io_br_taken_T) != $signed(_io_br_taken_T_1) : _GEN_264; // @[Decode.scala 557:23 Decode.scala 562:17]
  wire [63:0] _GEN_271 = 32'h1063 == _T_1 ? {{8'd0}, _io_br_target_T_5} : _GEN_265; // @[Decode.scala 557:23 Decode.scala 563:18]
  wire [5:0] _GEN_272 = 32'h4063 == _T_1 ? 6'h1 : _GEN_266; // @[Decode.scala 566:23 Decode.scala 567:15]
  wire  _GEN_273 = 32'h4063 == _T_1 | _GEN_267; // @[Decode.scala 566:23 Decode.scala 568:15]
  wire  _GEN_274 = 32'h4063 == _T_1 | _GEN_268; // @[Decode.scala 566:23 Decode.scala 569:15]
  wire  _GEN_275 = 32'h4063 == _T_1 ? 1'h0 : _GEN_269; // @[Decode.scala 566:23 Decode.scala 570:13]
  wire  _GEN_276 = 32'h4063 == _T_1 ? $signed(_io_br_taken_T) < $signed(_io_br_taken_T_1) : _GEN_270; // @[Decode.scala 566:23 Decode.scala 571:17]
  wire [63:0] _GEN_277 = 32'h4063 == _T_1 ? {{8'd0}, _io_br_target_T_5} : _GEN_271; // @[Decode.scala 566:23 Decode.scala 572:18]
  wire [5:0] _GEN_278 = 32'h5063 == _T_1 ? 6'h1 : _GEN_272; // @[Decode.scala 575:23 Decode.scala 576:15]
  wire  _GEN_279 = 32'h5063 == _T_1 | _GEN_273; // @[Decode.scala 575:23 Decode.scala 577:15]
  wire  _GEN_280 = 32'h5063 == _T_1 | _GEN_274; // @[Decode.scala 575:23 Decode.scala 578:15]
  wire  _GEN_281 = 32'h5063 == _T_1 ? 1'h0 : _GEN_275; // @[Decode.scala 575:23 Decode.scala 579:13]
  wire  _GEN_282 = 32'h5063 == _T_1 ? $signed(_io_br_taken_T) >= $signed(_io_br_taken_T_1) : _GEN_276; // @[Decode.scala 575:23 Decode.scala 580:17]
  wire [63:0] _GEN_283 = 32'h5063 == _T_1 ? {{8'd0}, _io_br_target_T_5} : _GEN_277; // @[Decode.scala 575:23 Decode.scala 581:18]
  wire [5:0] _GEN_284 = 32'h6063 == _T_1 ? 6'h1 : _GEN_278; // @[Decode.scala 584:24 Decode.scala 585:15]
  wire  _GEN_285 = 32'h6063 == _T_1 | _GEN_279; // @[Decode.scala 584:24 Decode.scala 586:15]
  wire  _GEN_286 = 32'h6063 == _T_1 | _GEN_280; // @[Decode.scala 584:24 Decode.scala 587:15]
  wire  _GEN_287 = 32'h6063 == _T_1 ? 1'h0 : _GEN_281; // @[Decode.scala 584:24 Decode.scala 588:13]
  wire  _GEN_288 = 32'h6063 == _T_1 ? rs1_value < rs2_value : _GEN_282; // @[Decode.scala 584:24 Decode.scala 589:17]
  wire [63:0] _GEN_289 = 32'h6063 == _T_1 ? {{8'd0}, _io_br_target_T_5} : _GEN_283; // @[Decode.scala 584:24 Decode.scala 590:18]
  wire [5:0] _GEN_290 = 32'h7063 == _T_1 ? 6'h1 : _GEN_284; // @[Decode.scala 593:24 Decode.scala 594:15]
  wire  _GEN_291 = 32'h7063 == _T_1 | _GEN_285; // @[Decode.scala 593:24 Decode.scala 595:15]
  wire  _GEN_292 = 32'h7063 == _T_1 | _GEN_286; // @[Decode.scala 593:24 Decode.scala 596:15]
  wire  _GEN_293 = 32'h7063 == _T_1 ? 1'h0 : _GEN_287; // @[Decode.scala 593:24 Decode.scala 597:13]
  wire [63:0] _GEN_295 = 32'h7063 == _T_1 ? {{8'd0}, _io_br_target_T_5} : _GEN_289; // @[Decode.scala 593:24 Decode.scala 599:18]
  wire  _T_114 = 32'h7b == id_inst; // @[Decode.scala 602:14]
  wire [5:0] id_opcode = 32'h7b == id_inst ? 6'h10 : _GEN_290; // @[Decode.scala 602:27 Decode.scala 605:15]
  wire [31:0] _id_op1_T_2 = _T_64 ? id_pc : 32'h0; // @[Decode.scala 624:31]
  wire [63:0] _id_op1_T_4 = 6'h10 == id_opcode ? rs1_value : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _id_op1_T_6 = 6'h20 == id_opcode ? {{32'd0}, _id_op1_T_2} : _id_op1_T_4; // @[Mux.scala 80:57]
  wire [63:0] _id_op1_T_8 = 6'h2 == id_opcode ? {{32'd0}, id_pc} : _id_op1_T_6; // @[Mux.scala 80:57]
  wire [63:0] _id_op1_T_10 = 6'h8 == id_opcode ? rs1_value : _id_op1_T_8; // @[Mux.scala 80:57]
  wire [63:0] _id_op1_T_12 = 6'h1 == id_opcode ? rs1_value : _id_op1_T_10; // @[Mux.scala 80:57]
  wire [63:0] id_op1 = 6'h4 == id_opcode ? rs1_value : _id_op1_T_12; // @[Mux.scala 80:57]
  wire  _GEN_301 = 32'h7b == id_inst ? 1'h0 : _GEN_293; // @[Decode.scala 602:27 Decode.scala 608:13]
  wire  id_wen = instr_valid & io_time_int ? 1'h0 : _GEN_301; // @[Decode.scala 611:37 Decode.scala 612:13]
  wire [3:0] id_sysop = instr_valid & io_time_int ? 4'h7 : _GEN_259; // @[Decode.scala 611:37 Decode.scala 613:14]
  wire  id_skip = _T_114 | id_inst == 32'h0; // @[Decode.scala 616:31]
  wire  _io_br_stall_T_11 = io_mem_stall & _rs2_forward_T & _rs2_forward_T_1 & io_rs2_en & id_valid_in; // @[Decode.scala 620:103]
  wire [63:0] _id_op2_T_1 = 6'h10 == id_opcode ? imm_i : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _id_op2_T_3 = 6'h20 == id_opcode ? imm_u : _id_op2_T_1; // @[Mux.scala 80:57]
  wire [63:0] _id_op2_T_5 = 6'h2 == id_opcode ? 64'h4 : _id_op2_T_3; // @[Mux.scala 80:57]
  wire [63:0] _id_op2_T_7 = 6'h8 == id_opcode ? rs2_value : _id_op2_T_5; // @[Mux.scala 80:57]
  wire [63:0] _id_op2_T_9 = 6'h1 == id_opcode ? rs2_value : _id_op2_T_7; // @[Mux.scala 80:57]
  assign io_rs1_addr = io_inst_my ? 5'ha : id_inst[19:15]; // @[Decode.scala 98:21]
  assign io_rs1_en = 32'h7b == id_inst | _GEN_291; // @[Decode.scala 602:27 Decode.scala 606:15]
  assign io_rs2_addr = id_inst[24:20]; // @[Decode.scala 99:22]
  assign io_rs2_en = 32'h7b == id_inst ? 1'h0 : _GEN_292; // @[Decode.scala 602:27 Decode.scala 607:15]
  assign io_id_pc = id_pc; // @[Decode.scala 641:15]
  assign io_id_inst = id_inst; // @[Decode.scala 642:15]
  assign io_id_wen = instr_valid & io_time_int ? 1'h0 : _GEN_301; // @[Decode.scala 611:37 Decode.scala 612:13]
  assign io_id_wdest = id_wen ? imm_s_lo : 5'h0; // @[Decode.scala 639:18]
  assign io_id_op1 = 6'h4 == id_opcode ? rs1_value : _id_op1_T_12; // @[Mux.scala 80:57]
  assign io_id_op2 = 6'h4 == id_opcode ? imm_s : _id_op2_T_9; // @[Mux.scala 80:57]
  assign io_rs2_value = rs2_forward ? _rs2_value_T_1 : io_rs2_data; // @[Decode.scala 115:22]
  assign io_type_w = 32'h4000503b == _T_21 | _GEN_247; // @[Decode.scala 530:24 Decode.scala 536:15]
  assign io_idop_aluop = io_flush ? 12'h0 : id_aluop; // @[Decode.scala 651:25]
  assign io_idop_loadop = io_flush ? 7'h0 : id_loadop; // @[Decode.scala 652:25]
  assign io_idop_storeop = io_flush ? 4'h0 : id_storeop; // @[Decode.scala 653:25]
  assign io_idop_sysop = io_flush ? 4'h0 : id_sysop; // @[Decode.scala 654:25]
  assign io_inst_my = 32'h7b == id_inst; // @[Decode.scala 602:14]
  assign io_skip = io_flush ? 1'h0 : id_skip; // @[Decode.scala 655:25]
  assign io_print = 32'h7b == id_inst ? id_op1 : 64'h0; // @[Decode.scala 602:27 Decode.scala 604:15 Decode.scala 106:14]
  assign io_br_valid = id_valid_in & ~io_br_stall; // @[Decode.scala 60:28]
  assign io_br_taken = 32'h7063 == _T_1 ? rs1_value >= rs2_value : _GEN_288; // @[Decode.scala 593:24 Decode.scala 598:17]
  assign io_br_target = _GEN_295[31:0];
  assign io_br_stall = io_mem_stall & _rs1_forward_T & _rs1_forward_T_1 & io_rs1_en & id_valid_in | _io_br_stall_T_11; // @[Decode.scala 619:116]
  assign io_if_allow_out = ~id_valid_in | io_id_valid_out & io_id_allow_out; // @[Decode.scala 62:29]
  assign io_id_valid_out = id_valid_in & ~io_br_stall; // @[Decode.scala 60:28]
  always @(posedge clock) begin
    if (reset) begin // @[Decode.scala 52:28]
      id_valid_in <= 1'h0; // @[Decode.scala 52:28]
    end else if (id_allow_in) begin // @[Decode.scala 56:22]
      id_valid_in <= io_if_valid_out; // @[Decode.scala 57:17]
    end
    if (reset) begin // @[Decode.scala 65:25]
      id_pc <= 32'h0; // @[Decode.scala 65:25]
    end else if (id_allow_in & io_if_valid_out) begin // @[Decode.scala 75:40]
      if (io_flush) begin // @[Decode.scala 76:19]
        id_pc <= 32'h0;
      end else begin
        id_pc <= io_fe_pc;
      end
    end
    if (reset) begin // @[Decode.scala 66:25]
      id_inst <= 32'h0; // @[Decode.scala 66:25]
    end else if (id_allow_in & io_if_valid_out) begin // @[Decode.scala 75:40]
      if (io_flush) begin // @[Decode.scala 77:19]
        id_inst <= 32'h0;
      end else begin
        id_inst <= io_fe_inst;
      end
    end
    if (reset) begin // @[Decode.scala 71:28]
      instr_valid <= 1'h0; // @[Decode.scala 71:28]
    end else if (id_allow_in & io_if_valid_out) begin // @[Decode.scala 75:40]
      instr_valid <= io_instr_valid; // @[Decode.scala 78:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  id_valid_in = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  id_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  id_inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  instr_valid = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Execution(
  input         clock,
  input         reset,
  input         io_type_w,
  input  [63:0] io_csr_rdata,
  input  [11:0] io_idop_aluop,
  input  [6:0]  io_idop_loadop,
  input  [3:0]  io_idop_storeop,
  input  [3:0]  io_idop_sysop,
  input  [31:0] io_id_pc,
  input  [31:0] io_id_inst,
  input         io_id_wen,
  input  [4:0]  io_id_wdest,
  input  [63:0] io_id_op1,
  input  [63:0] io_id_op2,
  output [31:0] io_ex_pc,
  output [31:0] io_ex_inst,
  output        io_ex_wen,
  output [4:0]  io_ex_wdest,
  output [63:0] io_ex_wdata,
  output [63:0] io_ex_op1,
  output        io_dmem_data_valid,
  input         io_dmem_data_ready,
  output        io_dmem_data_req,
  output [31:0] io_dmem_data_addr,
  output [1:0]  io_dmem_data_size,
  output [7:0]  io_dmem_data_strb,
  input  [63:0] io_dmem_data_read,
  output [63:0] io_dmem_data_write,
  input  [63:0] io_rs2_value,
  output [3:0]  io_ex_sysop,
  input         io_id_skip,
  output        io_cmp_ren,
  output        io_cmp_wen,
  output [63:0] io_cmp_addr,
  output [63:0] io_cmp_wdata,
  input  [63:0] io_cmp_rdata,
  input         io_flush,
  output        io_skip,
  output        io_mem_stall,
  output [4:0]  io_EX_wdest,
  output [63:0] io_EX_result,
  output        io_id_allow_out,
  output        io_ex_valid_out,
  input         io_id_valid_out,
  input         io_ex_allow_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg  ex_valid_in; // @[Execution.scala 51:28]
  reg  type_w; // @[Execution.scala 84:25]
  reg [11:0] ex_aluop; // @[Execution.scala 86:28]
  reg [63:0] ex_op1; // @[Execution.scala 81:25]
  wire [31:0] in1_hi = ex_op1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] in1_lo = ex_op1[31:0]; // @[Execution.scala 113:90]
  wire [63:0] _in1_T_3 = {in1_hi,in1_lo}; // @[Cat.scala 30:58]
  wire [63:0] _in1_T_4 = {32'h0,in1_lo}; // @[Cat.scala 30:58]
  wire [63:0] _in1_T_5 = ex_aluop == 12'h200 ? _in1_T_3 : _in1_T_4; // @[Execution.scala 113:28]
  wire [63:0] in1 = type_w ? _in1_T_5 : ex_op1; // @[Execution.scala 113:16]
  wire [63:0] _alu_result_0_T_14 = type_w ? _in1_T_5 : ex_op1; // @[Execution.scala 128:35]
  reg [63:0] ex_op2; // @[Execution.scala 82:25]
  wire [5:0] shamt = type_w ? {{1'd0}, ex_op2[4:0]} : ex_op2[5:0]; // @[Execution.scala 116:15]
  wire [63:0] _alu_result_0_T_16 = $signed(_alu_result_0_T_14) >>> shamt; // @[Execution.scala 128:54]
  wire [63:0] _alu_result_0_T_13 = in1 >> shamt; // @[Execution.scala 127:29]
  wire [126:0] _GEN_16 = {{63'd0}, in1}; // @[Execution.scala 126:30]
  wire [126:0] _alu_result_0_T_11 = _GEN_16 << shamt; // @[Execution.scala 126:30]
  wire [63:0] _alu_result_0_T_10 = in1 & ex_op2; // @[Execution.scala 125:29]
  wire [63:0] _alu_result_0_T_9 = in1 | ex_op2; // @[Execution.scala 124:29]
  wire [63:0] _alu_result_0_T_8 = in1 ^ ex_op2; // @[Execution.scala 123:29]
  wire  _alu_result_0_T_7 = in1 < ex_op2; // @[Execution.scala 122:29]
  wire  _alu_result_0_T_6 = $signed(_alu_result_0_T_14) < $signed(ex_op2); // @[Execution.scala 121:38]
  wire [63:0] _alu_result_0_T_3 = in1 - ex_op2; // @[Execution.scala 120:29]
  wire [63:0] _alu_result_0_T_1 = in1 + ex_op2; // @[Execution.scala 119:29]
  wire [63:0] _alu_result_0_T_18 = 12'h1 == ex_aluop ? _alu_result_0_T_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_20 = 12'h2 == ex_aluop ? _alu_result_0_T_3 : _alu_result_0_T_18; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_22 = 12'h4 == ex_aluop ? {{63'd0}, _alu_result_0_T_6} : _alu_result_0_T_20; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_24 = 12'h8 == ex_aluop ? {{63'd0}, _alu_result_0_T_7} : _alu_result_0_T_22; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_26 = 12'h10 == ex_aluop ? _alu_result_0_T_8 : _alu_result_0_T_24; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_28 = 12'h20 == ex_aluop ? _alu_result_0_T_9 : _alu_result_0_T_26; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_30 = 12'h40 == ex_aluop ? _alu_result_0_T_10 : _alu_result_0_T_28; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_32 = 12'h80 == ex_aluop ? _alu_result_0_T_11[63:0] : _alu_result_0_T_30; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_34 = 12'h100 == ex_aluop ? _alu_result_0_T_13 : _alu_result_0_T_32; // @[Mux.scala 80:57]
  wire [63:0] alu_result_0 = 12'h200 == ex_aluop ? _alu_result_0_T_16 : _alu_result_0_T_34; // @[Mux.scala 80:57]
  wire [31:0] alu_result_hi = alu_result_0[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] alu_result_lo = alu_result_0[31:0]; // @[Execution.scala 130:73]
  wire [63:0] _alu_result_T_2 = {alu_result_hi,alu_result_lo}; // @[Cat.scala 30:58]
  wire [63:0] alu_result = type_w ? _alu_result_T_2 : alu_result_0; // @[Execution.scala 130:20]
  wire [31:0] cmp_addr = alu_result[31:0];
  wire  _cmp_ren_T_2 = cmp_addr == 32'h2004000 | cmp_addr == 32'h200bff8; // @[Execution.scala 56:61]
  reg [6:0] ex_loadop; // @[Execution.scala 87:28]
  wire  load_en = ex_loadop != 7'h0; // @[Execution.scala 209:26]
  wire  cmp_ren = load_en & (cmp_addr == 32'h2004000 | cmp_addr == 32'h200bff8); // @[Execution.scala 56:28]
  reg [3:0] ex_storeop; // @[Execution.scala 88:28]
  wire  store_en = ex_storeop != 4'h0; // @[Execution.scala 210:27]
  wire  cmp_wen = store_en & _cmp_ren_T_2; // @[Execution.scala 57:28]
  wire  ex_allow_in = ~ex_valid_in | io_ex_valid_out & io_ex_allow_out; // @[Execution.scala 73:29]
  reg [31:0] ex_pc; // @[Execution.scala 76:25]
  reg [31:0] ex_inst; // @[Execution.scala 77:25]
  reg  ex_wen; // @[Execution.scala 78:25]
  reg [4:0] ex_wdest; // @[Execution.scala 79:25]
  reg [63:0] rs2_value; // @[Execution.scala 83:25]
  reg [3:0] ex_sysop; // @[Execution.scala 89:28]
  reg  ex_skip; // @[Execution.scala 90:28]
  wire [63:0] data_read = cmp_ren ? io_cmp_rdata : io_dmem_data_read; // @[Execution.scala 227:20]
  wire [55:0] mem_wdata_lb_hi = data_read[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mem_wdata_lb_lo = data_read[7:0]; // @[Execution.scala 140:56]
  wire [63:0] mem_wdata_lb = {mem_wdata_lb_hi,mem_wdata_lb_lo}; // @[Cat.scala 30:58]
  wire [63:0] mem_wdata_lbu = {56'h0,mem_wdata_lb_lo}; // @[Cat.scala 30:58]
  wire [47:0] mem_wdata_lh_hi = data_read[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [15:0] mem_wdata_lh_lo = data_read[15:0]; // @[Execution.scala 142:56]
  wire [63:0] mem_wdata_lh = {mem_wdata_lh_hi,mem_wdata_lh_lo}; // @[Cat.scala 30:58]
  wire [63:0] mem_wdata_lhu = {48'h0,mem_wdata_lh_lo}; // @[Cat.scala 30:58]
  wire [31:0] mem_wdata_lw_hi = data_read[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] mem_wdata_lw_lo = data_read[31:0]; // @[Execution.scala 144:56]
  wire [63:0] mem_wdata_lw = {mem_wdata_lw_hi,mem_wdata_lw_lo}; // @[Cat.scala 30:58]
  wire [63:0] mem_wdata_lwu = {32'h0,mem_wdata_lw_lo}; // @[Cat.scala 30:58]
  wire [31:0] _mem_wdata_T = ex_inst & 32'h707f; // @[Execution.scala 147:34]
  wire  _mem_wdata_T_1 = 32'h3 == _mem_wdata_T; // @[Execution.scala 147:34]
  wire [63:0] _mem_wdata_T_3 = _mem_wdata_T_1 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_4 = _mem_wdata_T_3 & mem_wdata_lb; // @[Execution.scala 147:43]
  wire  _mem_wdata_T_6 = 32'h4003 == _mem_wdata_T; // @[Execution.scala 148:34]
  wire [63:0] _mem_wdata_T_8 = _mem_wdata_T_6 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_9 = _mem_wdata_T_8 & mem_wdata_lbu; // @[Execution.scala 148:43]
  wire [63:0] _mem_wdata_T_10 = _mem_wdata_T_4 | _mem_wdata_T_9; // @[Execution.scala 147:60]
  wire  _mem_wdata_T_12 = 32'h1003 == _mem_wdata_T; // @[Execution.scala 149:34]
  wire [63:0] _mem_wdata_T_14 = _mem_wdata_T_12 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_15 = _mem_wdata_T_14 & mem_wdata_lh; // @[Execution.scala 149:43]
  wire [63:0] _mem_wdata_T_16 = _mem_wdata_T_10 | _mem_wdata_T_15; // @[Execution.scala 148:60]
  wire  _mem_wdata_T_18 = 32'h5003 == _mem_wdata_T; // @[Execution.scala 150:34]
  wire [63:0] _mem_wdata_T_20 = _mem_wdata_T_18 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_21 = _mem_wdata_T_20 & mem_wdata_lhu; // @[Execution.scala 150:43]
  wire [63:0] _mem_wdata_T_22 = _mem_wdata_T_16 | _mem_wdata_T_21; // @[Execution.scala 149:60]
  wire  _mem_wdata_T_24 = 32'h2003 == _mem_wdata_T; // @[Execution.scala 151:34]
  wire [63:0] _mem_wdata_T_26 = _mem_wdata_T_24 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_27 = _mem_wdata_T_26 & mem_wdata_lw; // @[Execution.scala 151:43]
  wire [63:0] _mem_wdata_T_28 = _mem_wdata_T_22 | _mem_wdata_T_27; // @[Execution.scala 150:60]
  wire  _mem_wdata_T_30 = 32'h6003 == _mem_wdata_T; // @[Execution.scala 152:34]
  wire [63:0] _mem_wdata_T_32 = _mem_wdata_T_30 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_33 = _mem_wdata_T_32 & mem_wdata_lwu; // @[Execution.scala 152:43]
  wire [63:0] _mem_wdata_T_34 = _mem_wdata_T_28 | _mem_wdata_T_33; // @[Execution.scala 151:60]
  wire  _mem_wdata_T_36 = 32'h3003 == _mem_wdata_T; // @[Execution.scala 153:34]
  wire [63:0] _mem_wdata_T_38 = _mem_wdata_T_36 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_39 = _mem_wdata_T_38 & data_read; // @[Execution.scala 153:43]
  wire [63:0] mem_wdata = _mem_wdata_T_34 | _mem_wdata_T_39; // @[Execution.scala 152:60]
  wire [7:0] data_write_sb_lo = rs2_value[7:0]; // @[Execution.scala 165:45]
  wire [63:0] _data_write_sb_T_1 = {56'h0,data_write_sb_lo}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_2 = {48'h0,data_write_sb_lo,8'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_3 = {40'h0,data_write_sb_lo,16'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_4 = {32'h0,data_write_sb_lo,24'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_5 = {24'h0,data_write_sb_lo,32'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_6 = {16'h0,data_write_sb_lo,40'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_7 = {8'h0,data_write_sb_lo,48'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_8 = {data_write_sb_lo,56'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_10 = 3'h1 == alu_result[2:0] ? _data_write_sb_T_2 : _data_write_sb_T_1; // @[Mux.scala 80:57]
  wire [63:0] _data_write_sb_T_12 = 3'h2 == alu_result[2:0] ? _data_write_sb_T_3 : _data_write_sb_T_10; // @[Mux.scala 80:57]
  wire [63:0] _data_write_sb_T_14 = 3'h3 == alu_result[2:0] ? _data_write_sb_T_4 : _data_write_sb_T_12; // @[Mux.scala 80:57]
  wire [63:0] _data_write_sb_T_16 = 3'h4 == alu_result[2:0] ? _data_write_sb_T_5 : _data_write_sb_T_14; // @[Mux.scala 80:57]
  wire [63:0] _data_write_sb_T_18 = 3'h5 == alu_result[2:0] ? _data_write_sb_T_6 : _data_write_sb_T_16; // @[Mux.scala 80:57]
  wire [63:0] _data_write_sb_T_20 = 3'h6 == alu_result[2:0] ? _data_write_sb_T_7 : _data_write_sb_T_18; // @[Mux.scala 80:57]
  wire [63:0] data_write_sb = 3'h7 == alu_result[2:0] ? _data_write_sb_T_8 : _data_write_sb_T_20; // @[Mux.scala 80:57]
  wire [1:0] _data_strb_sb_T_2 = 3'h1 == alu_result[2:0] ? 2'h2 : 2'h1; // @[Mux.scala 80:57]
  wire [2:0] _data_strb_sb_T_4 = 3'h2 == alu_result[2:0] ? 3'h4 : {{1'd0}, _data_strb_sb_T_2}; // @[Mux.scala 80:57]
  wire [3:0] _data_strb_sb_T_6 = 3'h3 == alu_result[2:0] ? 4'h8 : {{1'd0}, _data_strb_sb_T_4}; // @[Mux.scala 80:57]
  wire [4:0] _data_strb_sb_T_8 = 3'h4 == alu_result[2:0] ? 5'h10 : {{1'd0}, _data_strb_sb_T_6}; // @[Mux.scala 80:57]
  wire [5:0] _data_strb_sb_T_10 = 3'h5 == alu_result[2:0] ? 6'h20 : {{1'd0}, _data_strb_sb_T_8}; // @[Mux.scala 80:57]
  wire [6:0] _data_strb_sb_T_12 = 3'h6 == alu_result[2:0] ? 7'h40 : {{1'd0}, _data_strb_sb_T_10}; // @[Mux.scala 80:57]
  wire [7:0] data_strb_sb = 3'h7 == alu_result[2:0] ? 8'h80 : {{1'd0}, _data_strb_sb_T_12}; // @[Mux.scala 80:57]
  wire [15:0] data_write_sh_lo = rs2_value[15:0]; // @[Execution.scala 186:44]
  wire [63:0] _data_write_sh_T_1 = {48'h0,data_write_sh_lo}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sh_T_2 = {32'h0,data_write_sh_lo,16'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sh_T_3 = {16'h0,data_write_sh_lo,32'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sh_T_4 = {data_write_sh_lo,48'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sh_T_6 = 2'h1 == alu_result[2:1] ? _data_write_sh_T_2 : _data_write_sh_T_1; // @[Mux.scala 80:57]
  wire [63:0] _data_write_sh_T_8 = 2'h2 == alu_result[2:1] ? _data_write_sh_T_3 : _data_write_sh_T_6; // @[Mux.scala 80:57]
  wire [63:0] data_write_sh = 2'h3 == alu_result[2:1] ? _data_write_sh_T_4 : _data_write_sh_T_8; // @[Mux.scala 80:57]
  wire [3:0] _data_strb_sh_T_2 = 2'h1 == alu_result[2:1] ? 4'hc : 4'h3; // @[Mux.scala 80:57]
  wire [5:0] _data_strb_sh_T_4 = 2'h2 == alu_result[2:1] ? 6'h30 : {{2'd0}, _data_strb_sh_T_2}; // @[Mux.scala 80:57]
  wire [7:0] data_strb_sh = 2'h3 == alu_result[2:1] ? 8'hc0 : {{2'd0}, _data_strb_sh_T_4}; // @[Mux.scala 80:57]
  wire [32:0] data_write_sw_lo = rs2_value[32:0]; // @[Execution.scala 199:43]
  wire [64:0] _data_write_sw_T_1 = {32'h0,data_write_sw_lo}; // @[Cat.scala 30:58]
  wire [64:0] _data_write_sw_T_2 = {data_write_sw_lo,32'h0}; // @[Cat.scala 30:58]
  wire [64:0] _data_write_sw_T_4 = alu_result[2] ? _data_write_sw_T_2 : _data_write_sw_T_1; // @[Mux.scala 80:57]
  wire [7:0] data_strb_sw = alu_result[2] ? 8'hf0 : 8'hf; // @[Mux.scala 80:57]
  wire  _data_valid_T = load_en | store_en; // @[Execution.scala 212:26]
  wire  _data_write_T_1 = 32'h3023 == _mem_wdata_T; // @[Execution.scala 215:35]
  wire [63:0] _data_write_T_3 = _data_write_T_1 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _data_write_T_4 = _data_write_T_3 & rs2_value; // @[Execution.scala 215:43]
  wire  _data_write_T_6 = 32'h2023 == _mem_wdata_T; // @[Execution.scala 216:35]
  wire [63:0] _data_write_T_8 = _data_write_T_6 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] data_write_sw = _data_write_sw_T_4[63:0]; // @[Execution.scala 158:27 Execution.scala 198:17]
  wire [63:0] _data_write_T_9 = _data_write_T_8 & data_write_sw; // @[Execution.scala 216:43]
  wire [63:0] _data_write_T_10 = _data_write_T_4 | _data_write_T_9; // @[Execution.scala 215:60]
  wire  _data_write_T_12 = 32'h1023 == _mem_wdata_T; // @[Execution.scala 217:35]
  wire [63:0] _data_write_T_14 = _data_write_T_12 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _data_write_T_15 = _data_write_T_14 & data_write_sh; // @[Execution.scala 217:43]
  wire [63:0] _data_write_T_16 = _data_write_T_10 | _data_write_T_15; // @[Execution.scala 216:60]
  wire  _data_write_T_18 = 32'h23 == _mem_wdata_T; // @[Execution.scala 218:35]
  wire [63:0] _data_write_T_20 = _data_write_T_18 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _data_write_T_21 = _data_write_T_20 & data_write_sb; // @[Execution.scala 218:43]
  wire  _data_size_T_4 = _data_write_T_1 | _mem_wdata_T_36; // @[Execution.scala 219:42]
  wire [1:0] _data_size_T_6 = _data_size_T_4 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _data_size_T_15 = _data_write_T_6 | _mem_wdata_T_24 | _mem_wdata_T_30; // @[Execution.scala 220:60]
  wire [1:0] _data_size_T_17 = _data_size_T_15 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _data_size_T_18 = _data_size_T_17 & 2'h2; // @[Execution.scala 220:80]
  wire [1:0] _data_size_T_19 = _data_size_T_6 | _data_size_T_18; // @[Execution.scala 219:71]
  wire  _data_size_T_27 = _data_write_T_12 | _mem_wdata_T_12 | _mem_wdata_T_18; // @[Execution.scala 221:60]
  wire [1:0] _data_size_T_29 = _data_size_T_27 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _data_size_T_30 = _data_size_T_29 & 2'h1; // @[Execution.scala 221:80]
  wire [7:0] _data_strb_T_3 = _data_write_T_1 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _data_strb_T_8 = _data_write_T_6 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _data_strb_T_9 = _data_strb_T_8 & data_strb_sw; // @[Execution.scala 224:43]
  wire [7:0] _data_strb_T_10 = _data_strb_T_3 | _data_strb_T_9; // @[Execution.scala 223:59]
  wire [7:0] _data_strb_T_14 = _data_write_T_12 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _data_strb_T_15 = _data_strb_T_14 & data_strb_sh; // @[Execution.scala 225:43]
  wire [7:0] _data_strb_T_16 = _data_strb_T_10 | _data_strb_T_15; // @[Execution.scala 224:59]
  wire [7:0] _data_strb_T_20 = _data_write_T_18 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _data_strb_T_21 = _data_strb_T_20 & data_strb_sb; // @[Execution.scala 226:43]
  wire [63:0] _io_ex_wdata_T_1 = ex_sysop != 4'h0 ? io_csr_rdata : alu_result; // @[Execution.scala 242:45]
  assign io_ex_pc = io_flush ? 32'h0 : ex_pc; // @[Execution.scala 238:21]
  assign io_ex_inst = io_flush ? 32'h0 : ex_inst; // @[Execution.scala 239:21]
  assign io_ex_wen = io_flush ? 1'h0 : ex_wen; // @[Execution.scala 240:21]
  assign io_ex_wdest = ex_wdest; // @[Execution.scala 241:15]
  assign io_ex_wdata = load_en ? mem_wdata : _io_ex_wdata_T_1; // @[Execution.scala 242:21]
  assign io_ex_op1 = ex_op1; // @[Execution.scala 243:15]
  assign io_dmem_data_valid = (load_en | store_en) & (ex_valid_in & io_ex_allow_out) & (~cmp_ren & ~cmp_wen); // @[Execution.scala 212:72]
  assign io_dmem_data_req = ex_storeop != 4'h0; // @[Execution.scala 210:27]
  assign io_dmem_data_addr = alu_result[31:0]; // @[Execution.scala 232:23]
  assign io_dmem_data_size = _data_size_T_19 | _data_size_T_30; // @[Execution.scala 220:90]
  assign io_dmem_data_strb = _data_strb_T_16 | _data_strb_T_21; // @[Execution.scala 225:59]
  assign io_dmem_data_write = _data_write_T_16 | _data_write_T_21; // @[Execution.scala 217:60]
  assign io_ex_sysop = io_flush ? 4'h0 : ex_sysop; // @[Execution.scala 245:21]
  assign io_cmp_ren = load_en & (cmp_addr == 32'h2004000 | cmp_addr == 32'h200bff8); // @[Execution.scala 56:28]
  assign io_cmp_wen = store_en & _cmp_ren_T_2; // @[Execution.scala 57:28]
  assign io_cmp_addr = {{32'd0}, cmp_addr}; // @[Execution.scala 63:17]
  assign io_cmp_wdata = _data_write_T_16 | _data_write_T_21; // @[Execution.scala 217:60]
  assign io_skip = ex_skip | cmp_ren | cmp_wen; // @[Execution.scala 110:37]
  assign io_mem_stall = _data_valid_T & ~io_dmem_data_ready; // @[Execution.scala 250:41]
  assign io_EX_wdest = ex_valid_in ? ex_wdest : 5'h0; // @[Execution.scala 247:22]
  assign io_EX_result = io_ex_wdata; // @[Execution.scala 248:16]
  assign io_id_allow_out = ~ex_valid_in | io_ex_valid_out & io_ex_allow_out; // @[Execution.scala 73:29]
  assign io_ex_valid_out = ex_valid_in & (~load_en & ~store_en | io_dmem_data_ready | cmp_ren | cmp_wen | io_flush); // @[Execution.scala 71:28]
  always @(posedge clock) begin
    if (reset) begin // @[Execution.scala 51:28]
      ex_valid_in <= 1'h0; // @[Execution.scala 51:28]
    end else if (ex_allow_in) begin // @[Execution.scala 67:22]
      ex_valid_in <= io_id_valid_out; // @[Execution.scala 68:17]
    end
    if (reset) begin // @[Execution.scala 84:25]
      type_w <= 1'h0; // @[Execution.scala 84:25]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      type_w <= io_type_w; // @[Execution.scala 101:15]
    end
    if (reset) begin // @[Execution.scala 86:28]
      ex_aluop <= 12'h0; // @[Execution.scala 86:28]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      ex_aluop <= io_idop_aluop; // @[Execution.scala 103:15]
    end
    if (reset) begin // @[Execution.scala 81:25]
      ex_op1 <= 64'h0; // @[Execution.scala 81:25]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      ex_op1 <= io_id_op1; // @[Execution.scala 98:15]
    end
    if (reset) begin // @[Execution.scala 82:25]
      ex_op2 <= 64'h0; // @[Execution.scala 82:25]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      ex_op2 <= io_id_op2; // @[Execution.scala 99:15]
    end
    if (reset) begin // @[Execution.scala 87:28]
      ex_loadop <= 7'h0; // @[Execution.scala 87:28]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      ex_loadop <= io_idop_loadop; // @[Execution.scala 104:15]
    end
    if (reset) begin // @[Execution.scala 88:28]
      ex_storeop <= 4'h0; // @[Execution.scala 88:28]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      ex_storeop <= io_idop_storeop; // @[Execution.scala 105:15]
    end
    if (reset) begin // @[Execution.scala 76:25]
      ex_pc <= 32'h0; // @[Execution.scala 76:25]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      ex_pc <= io_id_pc; // @[Execution.scala 93:15]
    end
    if (reset) begin // @[Execution.scala 77:25]
      ex_inst <= 32'h0; // @[Execution.scala 77:25]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      ex_inst <= io_id_inst; // @[Execution.scala 94:15]
    end
    if (reset) begin // @[Execution.scala 78:25]
      ex_wen <= 1'h0; // @[Execution.scala 78:25]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      ex_wen <= io_id_wen; // @[Execution.scala 95:15]
    end
    if (reset) begin // @[Execution.scala 79:25]
      ex_wdest <= 5'h0; // @[Execution.scala 79:25]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      ex_wdest <= io_id_wdest; // @[Execution.scala 96:15]
    end
    if (reset) begin // @[Execution.scala 83:25]
      rs2_value <= 64'h0; // @[Execution.scala 83:25]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      rs2_value <= io_rs2_value; // @[Execution.scala 100:15]
    end
    if (reset) begin // @[Execution.scala 89:28]
      ex_sysop <= 4'h0; // @[Execution.scala 89:28]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      ex_sysop <= io_idop_sysop; // @[Execution.scala 106:15]
    end
    if (reset) begin // @[Execution.scala 90:28]
      ex_skip <= 1'h0; // @[Execution.scala 90:28]
    end else if (ex_allow_in & io_id_valid_out) begin // @[Execution.scala 92:40]
      ex_skip <= io_id_skip; // @[Execution.scala 107:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ex_valid_in = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  type_w = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ex_aluop = _RAND_2[11:0];
  _RAND_3 = {2{`RANDOM}};
  ex_op1 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ex_op2 = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  ex_loadop = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  ex_storeop = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  ex_pc = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  ex_inst = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  ex_wen = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ex_wdest = _RAND_10[4:0];
  _RAND_11 = {2{`RANDOM}};
  rs2_value = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  ex_sysop = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  ex_skip = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WriteBack(
  input         clock,
  input         reset,
  input  [31:0] io_ex_pc,
  input  [31:0] io_ex_inst,
  input         io_ex_wen,
  input  [4:0]  io_ex_wdest,
  input  [63:0] io_ex_wdata,
  input  [63:0] io_ex_op1,
  output [31:0] io_wb_pc,
  output [31:0] io_wb_inst,
  output        io_wb_wen,
  output [4:0]  io_wb_wdest,
  output [63:0] io_wb_wdata,
  output [63:0] io_wb_op1,
  input  [3:0]  io_ex_sysop,
  output [3:0]  io_sysop,
  input         io_ex_skip,
  output        io_skip,
  output        io_flush,
  output        io_ready_cmt,
  output [4:0]  io_WB_wdest,
  output [63:0] io_WB_result,
  output        io_intr,
  output        io_ex_allow_out,
  input         io_ex_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  wb_valid_in; // @[WriteBack.scala 48:28]
  wire  wb_allow_in = ~wb_valid_in | wb_valid_in; // @[WriteBack.scala 57:29]
  reg [31:0] wb_pc; // @[WriteBack.scala 60:25]
  reg [31:0] wb_inst; // @[WriteBack.scala 61:25]
  reg  wb_wen; // @[WriteBack.scala 62:25]
  reg [4:0] wb_wdest; // @[WriteBack.scala 63:25]
  reg [63:0] wb_wdata; // @[WriteBack.scala 64:25]
  reg [63:0] wb_op1; // @[WriteBack.scala 65:25]
  reg [3:0] wb_sysop; // @[WriteBack.scala 67:25]
  reg  wb_skip; // @[WriteBack.scala 68:25]
  wire  _io_intr_T = wb_sysop == 4'h7; // @[WriteBack.scala 70:23]
  wire  _io_wb_wen_T = wb_sysop != 4'h7; // @[WriteBack.scala 87:37]
  assign io_wb_pc = wb_pc; // @[WriteBack.scala 85:15]
  assign io_wb_inst = wb_inst; // @[WriteBack.scala 86:15]
  assign io_wb_wen = wb_wen & wb_sysop != 4'h7; // @[WriteBack.scala 87:25]
  assign io_wb_wdest = wb_wdest; // @[WriteBack.scala 88:15]
  assign io_wb_wdata = wb_wdata; // @[WriteBack.scala 89:15]
  assign io_wb_op1 = wb_op1; // @[WriteBack.scala 90:15]
  assign io_sysop = wb_sysop; // @[WriteBack.scala 92:15]
  assign io_skip = wb_skip; // @[WriteBack.scala 93:15]
  assign io_flush = (wb_sysop == 4'h4 | wb_sysop == 4'h5 | _io_intr_T) & wb_valid_in; // @[WriteBack.scala 95:110]
  assign io_ready_cmt = wb_valid_in & wb_inst != 32'h0 & _io_wb_wen_T; // @[WriteBack.scala 97:49]
  assign io_WB_wdest = wb_valid_in ? wb_wdest : 5'h0; // @[WriteBack.scala 99:22]
  assign io_WB_result = wb_wdata; // @[WriteBack.scala 100:16]
  assign io_intr = wb_sysop == 4'h7 & wb_valid_in; // @[WriteBack.scala 70:42]
  assign io_ex_allow_out = ~wb_valid_in | wb_valid_in; // @[WriteBack.scala 57:29]
  always @(posedge clock) begin
    if (reset) begin // @[WriteBack.scala 48:28]
      wb_valid_in <= 1'h0; // @[WriteBack.scala 48:28]
    end else if (wb_allow_in) begin // @[WriteBack.scala 52:22]
      wb_valid_in <= io_ex_valid_out; // @[WriteBack.scala 53:17]
    end
    if (reset) begin // @[WriteBack.scala 60:25]
      wb_pc <= 32'h0; // @[WriteBack.scala 60:25]
    end else if (wb_allow_in & io_ex_valid_out) begin // @[WriteBack.scala 73:40]
      wb_pc <= io_ex_pc; // @[WriteBack.scala 74:13]
    end
    if (reset) begin // @[WriteBack.scala 61:25]
      wb_inst <= 32'h0; // @[WriteBack.scala 61:25]
    end else if (wb_allow_in & io_ex_valid_out) begin // @[WriteBack.scala 73:40]
      wb_inst <= io_ex_inst; // @[WriteBack.scala 75:13]
    end
    if (reset) begin // @[WriteBack.scala 62:25]
      wb_wen <= 1'h0; // @[WriteBack.scala 62:25]
    end else if (wb_allow_in & io_ex_valid_out) begin // @[WriteBack.scala 73:40]
      wb_wen <= io_ex_wen; // @[WriteBack.scala 76:13]
    end
    if (reset) begin // @[WriteBack.scala 63:25]
      wb_wdest <= 5'h0; // @[WriteBack.scala 63:25]
    end else if (wb_allow_in & io_ex_valid_out) begin // @[WriteBack.scala 73:40]
      wb_wdest <= io_ex_wdest; // @[WriteBack.scala 77:13]
    end
    if (reset) begin // @[WriteBack.scala 64:25]
      wb_wdata <= 64'h0; // @[WriteBack.scala 64:25]
    end else if (wb_allow_in & io_ex_valid_out) begin // @[WriteBack.scala 73:40]
      wb_wdata <= io_ex_wdata; // @[WriteBack.scala 78:13]
    end
    if (reset) begin // @[WriteBack.scala 65:25]
      wb_op1 <= 64'h0; // @[WriteBack.scala 65:25]
    end else if (wb_allow_in & io_ex_valid_out) begin // @[WriteBack.scala 73:40]
      wb_op1 <= io_ex_op1; // @[WriteBack.scala 79:13]
    end
    if (reset) begin // @[WriteBack.scala 67:25]
      wb_sysop <= 4'h0; // @[WriteBack.scala 67:25]
    end else if (wb_allow_in & io_ex_valid_out) begin // @[WriteBack.scala 73:40]
      wb_sysop <= io_ex_sysop; // @[WriteBack.scala 81:13]
    end
    if (reset) begin // @[WriteBack.scala 68:25]
      wb_skip <= 1'h0; // @[WriteBack.scala 68:25]
    end else if (wb_allow_in & io_ex_valid_out) begin // @[WriteBack.scala 73:40]
      wb_skip <= io_ex_skip; // @[WriteBack.scala 82:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wb_valid_in = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wb_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  wb_inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  wb_wen = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wb_wdest = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  wb_wdata = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  wb_op1 = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  wb_sysop = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  wb_skip = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_rs1_addr,
  input  [4:0]  io_rs2_addr,
  output [63:0] io_rs1_data,
  output [63:0] io_rs2_data,
  input  [4:0]  io_rd_addr,
  input  [63:0] io_rd_data,
  input         io_rd_en,
  output [63:0] rf_10
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire  dt_ar_clock; // @[RegFile.scala 25:21]
  wire [7:0] dt_ar_coreid; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_0; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_1; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_2; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_3; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_4; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_5; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_6; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_7; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_8; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_9; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_10; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_11; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_12; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_13; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_14; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_15; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_16; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_17; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_18; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_19; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_20; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_21; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_22; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_23; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_24; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_25; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_26; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_27; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_28; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_29; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_30; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_31; // @[RegFile.scala 25:21]
  reg [63:0] rf__0; // @[RegFile.scala 16:19]
  reg [63:0] rf__1; // @[RegFile.scala 16:19]
  reg [63:0] rf__2; // @[RegFile.scala 16:19]
  reg [63:0] rf__3; // @[RegFile.scala 16:19]
  reg [63:0] rf__4; // @[RegFile.scala 16:19]
  reg [63:0] rf__5; // @[RegFile.scala 16:19]
  reg [63:0] rf__6; // @[RegFile.scala 16:19]
  reg [63:0] rf__7; // @[RegFile.scala 16:19]
  reg [63:0] rf__8; // @[RegFile.scala 16:19]
  reg [63:0] rf__9; // @[RegFile.scala 16:19]
  reg [63:0] rf__10; // @[RegFile.scala 16:19]
  reg [63:0] rf__11; // @[RegFile.scala 16:19]
  reg [63:0] rf__12; // @[RegFile.scala 16:19]
  reg [63:0] rf__13; // @[RegFile.scala 16:19]
  reg [63:0] rf__14; // @[RegFile.scala 16:19]
  reg [63:0] rf__15; // @[RegFile.scala 16:19]
  reg [63:0] rf__16; // @[RegFile.scala 16:19]
  reg [63:0] rf__17; // @[RegFile.scala 16:19]
  reg [63:0] rf__18; // @[RegFile.scala 16:19]
  reg [63:0] rf__19; // @[RegFile.scala 16:19]
  reg [63:0] rf__20; // @[RegFile.scala 16:19]
  reg [63:0] rf__21; // @[RegFile.scala 16:19]
  reg [63:0] rf__22; // @[RegFile.scala 16:19]
  reg [63:0] rf__23; // @[RegFile.scala 16:19]
  reg [63:0] rf__24; // @[RegFile.scala 16:19]
  reg [63:0] rf__25; // @[RegFile.scala 16:19]
  reg [63:0] rf__26; // @[RegFile.scala 16:19]
  reg [63:0] rf__27; // @[RegFile.scala 16:19]
  reg [63:0] rf__28; // @[RegFile.scala 16:19]
  reg [63:0] rf__29; // @[RegFile.scala 16:19]
  reg [63:0] rf__30; // @[RegFile.scala 16:19]
  reg [63:0] rf__31; // @[RegFile.scala 16:19]
  wire [63:0] _GEN_65 = 5'h1 == io_rs1_addr ? rf__1 : rf__0; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_66 = 5'h2 == io_rs1_addr ? rf__2 : _GEN_65; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_67 = 5'h3 == io_rs1_addr ? rf__3 : _GEN_66; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_68 = 5'h4 == io_rs1_addr ? rf__4 : _GEN_67; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_69 = 5'h5 == io_rs1_addr ? rf__5 : _GEN_68; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_70 = 5'h6 == io_rs1_addr ? rf__6 : _GEN_69; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_71 = 5'h7 == io_rs1_addr ? rf__7 : _GEN_70; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_72 = 5'h8 == io_rs1_addr ? rf__8 : _GEN_71; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_73 = 5'h9 == io_rs1_addr ? rf__9 : _GEN_72; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_74 = 5'ha == io_rs1_addr ? rf__10 : _GEN_73; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_75 = 5'hb == io_rs1_addr ? rf__11 : _GEN_74; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_76 = 5'hc == io_rs1_addr ? rf__12 : _GEN_75; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_77 = 5'hd == io_rs1_addr ? rf__13 : _GEN_76; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_78 = 5'he == io_rs1_addr ? rf__14 : _GEN_77; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_79 = 5'hf == io_rs1_addr ? rf__15 : _GEN_78; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_80 = 5'h10 == io_rs1_addr ? rf__16 : _GEN_79; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_81 = 5'h11 == io_rs1_addr ? rf__17 : _GEN_80; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_82 = 5'h12 == io_rs1_addr ? rf__18 : _GEN_81; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_83 = 5'h13 == io_rs1_addr ? rf__19 : _GEN_82; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_84 = 5'h14 == io_rs1_addr ? rf__20 : _GEN_83; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_85 = 5'h15 == io_rs1_addr ? rf__21 : _GEN_84; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_86 = 5'h16 == io_rs1_addr ? rf__22 : _GEN_85; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_87 = 5'h17 == io_rs1_addr ? rf__23 : _GEN_86; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_88 = 5'h18 == io_rs1_addr ? rf__24 : _GEN_87; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_89 = 5'h19 == io_rs1_addr ? rf__25 : _GEN_88; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_90 = 5'h1a == io_rs1_addr ? rf__26 : _GEN_89; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_91 = 5'h1b == io_rs1_addr ? rf__27 : _GEN_90; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_92 = 5'h1c == io_rs1_addr ? rf__28 : _GEN_91; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_93 = 5'h1d == io_rs1_addr ? rf__29 : _GEN_92; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_94 = 5'h1e == io_rs1_addr ? rf__30 : _GEN_93; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_95 = 5'h1f == io_rs1_addr ? rf__31 : _GEN_94; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_97 = 5'h1 == io_rs2_addr ? rf__1 : rf__0; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_98 = 5'h2 == io_rs2_addr ? rf__2 : _GEN_97; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_99 = 5'h3 == io_rs2_addr ? rf__3 : _GEN_98; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_100 = 5'h4 == io_rs2_addr ? rf__4 : _GEN_99; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_101 = 5'h5 == io_rs2_addr ? rf__5 : _GEN_100; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_102 = 5'h6 == io_rs2_addr ? rf__6 : _GEN_101; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_103 = 5'h7 == io_rs2_addr ? rf__7 : _GEN_102; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_104 = 5'h8 == io_rs2_addr ? rf__8 : _GEN_103; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_105 = 5'h9 == io_rs2_addr ? rf__9 : _GEN_104; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_106 = 5'ha == io_rs2_addr ? rf__10 : _GEN_105; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_107 = 5'hb == io_rs2_addr ? rf__11 : _GEN_106; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_108 = 5'hc == io_rs2_addr ? rf__12 : _GEN_107; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_109 = 5'hd == io_rs2_addr ? rf__13 : _GEN_108; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_110 = 5'he == io_rs2_addr ? rf__14 : _GEN_109; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_111 = 5'hf == io_rs2_addr ? rf__15 : _GEN_110; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_112 = 5'h10 == io_rs2_addr ? rf__16 : _GEN_111; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_113 = 5'h11 == io_rs2_addr ? rf__17 : _GEN_112; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_114 = 5'h12 == io_rs2_addr ? rf__18 : _GEN_113; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_115 = 5'h13 == io_rs2_addr ? rf__19 : _GEN_114; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_116 = 5'h14 == io_rs2_addr ? rf__20 : _GEN_115; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_117 = 5'h15 == io_rs2_addr ? rf__21 : _GEN_116; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_118 = 5'h16 == io_rs2_addr ? rf__22 : _GEN_117; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_119 = 5'h17 == io_rs2_addr ? rf__23 : _GEN_118; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_120 = 5'h18 == io_rs2_addr ? rf__24 : _GEN_119; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_121 = 5'h19 == io_rs2_addr ? rf__25 : _GEN_120; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_122 = 5'h1a == io_rs2_addr ? rf__26 : _GEN_121; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_123 = 5'h1b == io_rs2_addr ? rf__27 : _GEN_122; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_124 = 5'h1c == io_rs2_addr ? rf__28 : _GEN_123; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_125 = 5'h1d == io_rs2_addr ? rf__29 : _GEN_124; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_126 = 5'h1e == io_rs2_addr ? rf__30 : _GEN_125; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_127 = 5'h1f == io_rs2_addr ? rf__31 : _GEN_126; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  DifftestArchIntRegState dt_ar ( // @[RegFile.scala 25:21]
    .clock(dt_ar_clock),
    .coreid(dt_ar_coreid),
    .gpr_0(dt_ar_gpr_0),
    .gpr_1(dt_ar_gpr_1),
    .gpr_2(dt_ar_gpr_2),
    .gpr_3(dt_ar_gpr_3),
    .gpr_4(dt_ar_gpr_4),
    .gpr_5(dt_ar_gpr_5),
    .gpr_6(dt_ar_gpr_6),
    .gpr_7(dt_ar_gpr_7),
    .gpr_8(dt_ar_gpr_8),
    .gpr_9(dt_ar_gpr_9),
    .gpr_10(dt_ar_gpr_10),
    .gpr_11(dt_ar_gpr_11),
    .gpr_12(dt_ar_gpr_12),
    .gpr_13(dt_ar_gpr_13),
    .gpr_14(dt_ar_gpr_14),
    .gpr_15(dt_ar_gpr_15),
    .gpr_16(dt_ar_gpr_16),
    .gpr_17(dt_ar_gpr_17),
    .gpr_18(dt_ar_gpr_18),
    .gpr_19(dt_ar_gpr_19),
    .gpr_20(dt_ar_gpr_20),
    .gpr_21(dt_ar_gpr_21),
    .gpr_22(dt_ar_gpr_22),
    .gpr_23(dt_ar_gpr_23),
    .gpr_24(dt_ar_gpr_24),
    .gpr_25(dt_ar_gpr_25),
    .gpr_26(dt_ar_gpr_26),
    .gpr_27(dt_ar_gpr_27),
    .gpr_28(dt_ar_gpr_28),
    .gpr_29(dt_ar_gpr_29),
    .gpr_30(dt_ar_gpr_30),
    .gpr_31(dt_ar_gpr_31)
  );
  assign io_rs1_data = io_rs1_addr != 5'h0 ? _GEN_95 : 64'h0; // @[RegFile.scala 22:21]
  assign io_rs2_data = io_rs2_addr != 5'h0 ? _GEN_127 : 64'h0; // @[RegFile.scala 23:21]
  assign rf_10 = rf__10;
  assign dt_ar_clock = clock; // @[RegFile.scala 26:19]
  assign dt_ar_coreid = 8'h0; // @[RegFile.scala 27:19]
  assign dt_ar_gpr_0 = rf__0; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_1 = rf__1; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_2 = rf__2; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_3 = rf__3; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_4 = rf__4; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_5 = rf__5; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_6 = rf__6; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_7 = rf__7; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_8 = rf__8; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_9 = rf__9; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_10 = rf__10; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_11 = rf__11; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_12 = rf__12; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_13 = rf__13; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_14 = rf__14; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_15 = rf__15; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_16 = rf__16; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_17 = rf__17; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_18 = rf__18; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_19 = rf__19; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_20 = rf__20; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_21 = rf__21; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_22 = rf__22; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_23 = rf__23; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_24 = rf__24; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_25 = rf__25; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_26 = rf__26; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_27 = rf__27; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_28 = rf__28; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_29 = rf__29; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_30 = rf__30; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_31 = rf__31; // @[RegFile.scala 28:19]
  always @(posedge clock) begin
    if (reset) begin // @[RegFile.scala 16:19]
      rf__0 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h0 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__0 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__1 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__1 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__2 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h2 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__2 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__3 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h3 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__3 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__4 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h4 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__4 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__5 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h5 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__5 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__6 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h6 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__6 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__7 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h7 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__7 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__8 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h8 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__8 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__9 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h9 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__9 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__10 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'ha == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__10 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__11 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'hb == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__11 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__12 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'hc == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__12 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__13 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'hd == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__13 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__14 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'he == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__14 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__15 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'hf == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__15 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__16 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h10 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__16 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__17 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h11 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__17 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__18 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h12 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__18 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__19 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h13 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__19 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__20 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h14 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__20 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__21 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h15 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__21 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__22 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h16 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__22 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__23 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h17 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__23 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__24 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h18 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__24 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__25 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h19 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__25 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__26 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1a == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__26 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__27 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1b == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__27 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__28 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1c == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__28 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__29 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1d == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__29 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__30 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1e == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__30 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__31 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1f == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__31 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rf__0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  rf__1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf__2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf__3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf__4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf__5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf__6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf__7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf__8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf__9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf__10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf__11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf__12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf__13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf__14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf__15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf__16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf__17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf__18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf__19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf__20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf__21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf__22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf__23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf__24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf__25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf__26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf__27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf__28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf__29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf__30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  rf__31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Csr(
  input         clock,
  input         reset,
  input  [63:0] io_in1,
  input  [31:0] io_pc,
  input  [31:0] io_inst,
  input  [3:0]  io_sysop,
  output [63:0] io_csr_rdata,
  output        io_csr_jmp,
  output [31:0] io_newpc,
  output [63:0] io_mstatus,
  output [63:0] io_mie,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  dt_cs_clock; // @[Csr.scala 151:21]
  wire [7:0] dt_cs_coreid; // @[Csr.scala 151:21]
  wire [1:0] dt_cs_priviledgeMode; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_mstatus; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_sstatus; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_mepc; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_sepc; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_mtval; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_stval; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_mtvec; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_stvec; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_mcause; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_scause; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_satp; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_mip; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_mie; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_mscratch; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_sscratch; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_mideleg; // @[Csr.scala 151:21]
  wire [63:0] dt_cs_medeleg; // @[Csr.scala 151:21]
  wire [4:0] in2_lo = io_inst[19:15]; // @[Csr.scala 24:39]
  wire [63:0] in2 = {59'h0,in2_lo}; // @[Cat.scala 30:58]
  wire  _csr_rw_T = io_sysop == 4'h1; // @[Csr.scala 26:23]
  wire  _csr_rw_T_1 = io_sysop == 4'h2; // @[Csr.scala 27:23]
  wire  _csr_rw_T_2 = io_sysop == 4'h1 | _csr_rw_T_1; // @[Csr.scala 26:46]
  wire  _csr_rw_T_4 = _csr_rw_T_2 | _csr_rw_T; // @[Csr.scala 27:46]
  wire  _csr_rw_T_5 = io_sysop == 4'h8; // @[Csr.scala 29:23]
  wire  _csr_rw_T_6 = _csr_rw_T_4 | _csr_rw_T_5; // @[Csr.scala 28:46]
  wire  _csr_rw_T_7 = io_sysop == 4'h9; // @[Csr.scala 30:23]
  wire  csr_rw = _csr_rw_T_6 | _csr_rw_T_7; // @[Csr.scala 29:46]
  reg [63:0] mstatus; // @[Csr.scala 40:26]
  reg [63:0] mie; // @[Csr.scala 41:26]
  reg [63:0] mtvec; // @[Csr.scala 43:26]
  reg [63:0] mscratch; // @[Csr.scala 44:26]
  reg [63:0] mepc; // @[Csr.scala 45:26]
  reg [63:0] mcause; // @[Csr.scala 46:26]
  reg [63:0] mcycle; // @[Csr.scala 47:26]
  wire  _T_1 = io_sysop == 4'h4 & io_flush; // @[Csr.scala 61:36]
  wire [50:0] mstatus_hi_hi_hi = mstatus[63:13]; // @[Csr.scala 64:27]
  wire [2:0] mstatus_hi_lo_hi = mstatus[10:8]; // @[Csr.scala 64:57]
  wire  mstatus_hi_lo_lo = mstatus[3]; // @[Csr.scala 64:72]
  wire [2:0] mstatus_lo_hi_hi = mstatus[6:4]; // @[Csr.scala 64:84]
  wire [2:0] mstatus_lo_lo = mstatus[2:0]; // @[Csr.scala 64:104]
  wire [63:0] _mstatus_T = {mstatus_hi_hi_hi,2'h3,mstatus_hi_lo_hi,mstatus_hi_lo_lo,mstatus_lo_hi_hi,1'h0,mstatus_lo_lo}
    ; // @[Cat.scala 30:58]
  wire [29:0] newpc_hi = mtvec[31:2]; // @[Csr.scala 66:23]
  wire [31:0] _newpc_T = {newpc_hi,2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_0 = io_sysop == 4'h4 & io_flush ? {{32'd0}, io_pc} : mepc; // @[Csr.scala 61:49 Csr.scala 62:10 Csr.scala 45:26]
  wire [63:0] _GEN_1 = io_sysop == 4'h4 & io_flush ? 64'hb : mcause; // @[Csr.scala 61:49 Csr.scala 63:12 Csr.scala 46:26]
  wire [63:0] _GEN_2 = io_sysop == 4'h4 & io_flush ? _mstatus_T : mstatus; // @[Csr.scala 61:49 Csr.scala 64:13 Csr.scala 40:26]
  wire [31:0] _GEN_4 = io_sysop == 4'h4 & io_flush ? _newpc_T : 32'h0; // @[Csr.scala 61:49 Csr.scala 66:11]
  wire  mstatus_lo_hi_lo = mstatus[7]; // @[Csr.scala 71:92]
  wire [63:0] _mstatus_T_1 = {mstatus_hi_hi_hi,2'h0,mstatus_hi_lo_hi,1'h1,mstatus_lo_hi_hi,mstatus_lo_hi_lo,
    mstatus_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_5 = io_sysop == 4'h5 & io_flush ? _mstatus_T_1 : _GEN_2; // @[Csr.scala 70:48 Csr.scala 71:13]
  wire  _GEN_6 = io_sysop == 4'h5 & io_flush | _T_1; // @[Csr.scala 70:48 Csr.scala 72:13]
  wire [31:0] _GEN_7 = io_sysop == 4'h5 & io_flush ? mepc[31:0] : _GEN_4; // @[Csr.scala 70:48 Csr.scala 73:11]
  wire [63:0] _GEN_8 = io_sysop == 4'h7 & io_flush ? {{32'd0}, io_pc} : _GEN_0; // @[Csr.scala 77:47 Csr.scala 78:10]
  wire [63:0] _GEN_9 = io_sysop == 4'h7 & io_flush ? 64'h8000000000000007 : _GEN_1; // @[Csr.scala 77:47 Csr.scala 79:12]
  wire [63:0] _GEN_10 = io_sysop == 4'h7 & io_flush ? _mstatus_T : _GEN_5; // @[Csr.scala 77:47 Csr.scala 80:13]
  wire [63:0] _mcycle_T_1 = mcycle + 64'h1; // @[Csr.scala 87:20]
  wire [11:0] addr = io_inst[31:20]; // @[Csr.scala 91:21]
  wire [63:0] _rdata_T_1 = 12'h300 == addr ? mstatus : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_3 = 12'h342 == addr ? mcause : _rdata_T_1; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_5 = 12'h304 == addr ? mie : _rdata_T_3; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_7 = 12'h305 == addr ? mtvec : _rdata_T_5; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_9 = 12'h340 == addr ? mscratch : _rdata_T_7; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_11 = 12'h341 == addr ? mepc : _rdata_T_9; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_13 = 12'h344 == addr ? 64'h0 : _rdata_T_11; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_15 = 12'hb00 == addr ? mcycle : _rdata_T_13; // @[Mux.scala 80:57]
  wire [63:0] rdata = 12'hb02 == addr ? 64'h0 : _rdata_T_15; // @[Mux.scala 80:57]
  wire [63:0] _wdata_T = rdata | io_in1; // @[Csr.scala 98:33]
  wire [63:0] _wdata_T_1 = ~io_in1; // @[Csr.scala 99:35]
  wire [63:0] _wdata_T_2 = rdata & _wdata_T_1; // @[Csr.scala 99:33]
  wire [63:0] _wdata_T_3 = rdata | in2; // @[Csr.scala 100:33]
  wire [63:0] _wdata_T_4 = ~in2; // @[Csr.scala 101:35]
  wire [63:0] _wdata_T_5 = rdata & _wdata_T_4; // @[Csr.scala 101:33]
  wire [63:0] _wdata_T_7 = 4'h1 == io_sysop ? io_in1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _wdata_T_9 = 4'h2 == io_sysop ? _wdata_T : _wdata_T_7; // @[Mux.scala 80:57]
  wire [63:0] _wdata_T_11 = 4'h3 == io_sysop ? _wdata_T_2 : _wdata_T_9; // @[Mux.scala 80:57]
  wire [63:0] _wdata_T_13 = 4'h8 == io_sysop ? _wdata_T_3 : _wdata_T_11; // @[Mux.scala 80:57]
  wire [63:0] wdata = 4'h9 == io_sysop ? _wdata_T_5 : _wdata_T_13; // @[Mux.scala 80:57]
  wire  mstatus_hi_3 = wdata[16] & wdata[15] | wdata[14] & wdata[13]; // @[Csr.scala 134:46]
  wire [62:0] mstatus_lo_3 = wdata[62:0]; // @[Csr.scala 134:79]
  wire [63:0] _mstatus_T_9 = {mstatus_hi_3,mstatus_lo_3}; // @[Cat.scala 30:58]
  DifftestCSRState dt_cs ( // @[Csr.scala 151:21]
    .clock(dt_cs_clock),
    .coreid(dt_cs_coreid),
    .priviledgeMode(dt_cs_priviledgeMode),
    .mstatus(dt_cs_mstatus),
    .sstatus(dt_cs_sstatus),
    .mepc(dt_cs_mepc),
    .sepc(dt_cs_sepc),
    .mtval(dt_cs_mtval),
    .stval(dt_cs_stval),
    .mtvec(dt_cs_mtvec),
    .stvec(dt_cs_stvec),
    .mcause(dt_cs_mcause),
    .scause(dt_cs_scause),
    .satp(dt_cs_satp),
    .mip(dt_cs_mip),
    .mie(dt_cs_mie),
    .mscratch(dt_cs_mscratch),
    .sscratch(dt_cs_sscratch),
    .mideleg(dt_cs_mideleg),
    .medeleg(dt_cs_medeleg)
  );
  assign io_csr_rdata = 12'hb02 == addr ? 64'h0 : _rdata_T_15; // @[Mux.scala 80:57]
  assign io_csr_jmp = io_sysop == 4'h7 & io_flush | _GEN_6; // @[Csr.scala 77:47 Csr.scala 81:13]
  assign io_newpc = io_sysop == 4'h7 & io_flush ? _newpc_T : _GEN_7; // @[Csr.scala 77:47 Csr.scala 82:11]
  assign io_mstatus = mstatus; // @[Csr.scala 146:14]
  assign io_mie = mie; // @[Csr.scala 147:10]
  assign dt_cs_clock = clock; // @[Csr.scala 152:27]
  assign dt_cs_coreid = 8'h0; // @[Csr.scala 153:27]
  assign dt_cs_priviledgeMode = 2'h3; // @[Csr.scala 154:27]
  assign dt_cs_mstatus = mstatus; // @[Csr.scala 155:27]
  assign dt_cs_sstatus = mstatus & 64'h80000003000de122; // @[Csr.scala 156:38]
  assign dt_cs_mepc = mepc; // @[Csr.scala 157:27]
  assign dt_cs_sepc = 64'h0; // @[Csr.scala 158:27]
  assign dt_cs_mtval = 64'h0; // @[Csr.scala 159:27]
  assign dt_cs_stval = 64'h0; // @[Csr.scala 160:27]
  assign dt_cs_mtvec = mtvec; // @[Csr.scala 161:27]
  assign dt_cs_stvec = 64'h0; // @[Csr.scala 162:27]
  assign dt_cs_mcause = mcause; // @[Csr.scala 163:27]
  assign dt_cs_scause = 64'h0; // @[Csr.scala 164:27]
  assign dt_cs_satp = 64'h0; // @[Csr.scala 165:27]
  assign dt_cs_mip = 64'h0; // @[Csr.scala 166:27]
  assign dt_cs_mie = mie; // @[Csr.scala 167:27]
  assign dt_cs_mscratch = mscratch; // @[Csr.scala 168:27]
  assign dt_cs_sscratch = 64'h0; // @[Csr.scala 169:27]
  assign dt_cs_mideleg = 64'h0; // @[Csr.scala 170:27]
  assign dt_cs_medeleg = 64'h0; // @[Csr.scala 171:27]
  always @(posedge clock) begin
    if (reset) begin // @[Csr.scala 40:26]
      mstatus <= 64'h1800; // @[Csr.scala 40:26]
    end else if (csr_rw) begin // @[Csr.scala 118:13]
      if (addr == 12'h300) begin // @[Csr.scala 131:33]
        mstatus <= _mstatus_T_9; // @[Csr.scala 134:15]
      end else begin
        mstatus <= _GEN_10;
      end
    end else begin
      mstatus <= _GEN_10;
    end
    if (reset) begin // @[Csr.scala 41:26]
      mie <= 64'h0; // @[Csr.scala 41:26]
    end else if (csr_rw) begin // @[Csr.scala 118:13]
      if (addr == 12'h304) begin // @[Csr.scala 136:29]
        if (4'h9 == io_sysop) begin // @[Mux.scala 80:57]
          mie <= _wdata_T_5;
        end else begin
          mie <= _wdata_T_13;
        end
      end
    end
    if (reset) begin // @[Csr.scala 43:26]
      mtvec <= 64'h0; // @[Csr.scala 43:26]
    end else if (csr_rw) begin // @[Csr.scala 118:13]
      if (addr == 12'h305) begin // @[Csr.scala 122:31]
        if (4'h9 == io_sysop) begin // @[Mux.scala 80:57]
          mtvec <= _wdata_T_5;
        end else begin
          mtvec <= _wdata_T_13;
        end
      end
    end
    if (reset) begin // @[Csr.scala 44:26]
      mscratch <= 64'h0; // @[Csr.scala 44:26]
    end else if (csr_rw) begin // @[Csr.scala 118:13]
      if (addr == 12'h340) begin // @[Csr.scala 139:34]
        if (4'h9 == io_sysop) begin // @[Mux.scala 80:57]
          mscratch <= _wdata_T_5;
        end else begin
          mscratch <= _wdata_T_13;
        end
      end
    end
    if (reset) begin // @[Csr.scala 45:26]
      mepc <= 64'h0; // @[Csr.scala 45:26]
    end else if (csr_rw) begin // @[Csr.scala 118:13]
      if (addr == 12'h341) begin // @[Csr.scala 125:30]
        if (4'h9 == io_sysop) begin // @[Mux.scala 80:57]
          mepc <= _wdata_T_5;
        end else begin
          mepc <= _wdata_T_13;
        end
      end else begin
        mepc <= _GEN_8;
      end
    end else begin
      mepc <= _GEN_8;
    end
    if (reset) begin // @[Csr.scala 46:26]
      mcause <= 64'h0; // @[Csr.scala 46:26]
    end else if (csr_rw) begin // @[Csr.scala 118:13]
      if (addr == 12'h342) begin // @[Csr.scala 128:32]
        if (4'h9 == io_sysop) begin // @[Mux.scala 80:57]
          mcause <= _wdata_T_5;
        end else begin
          mcause <= _wdata_T_13;
        end
      end else begin
        mcause <= _GEN_9;
      end
    end else begin
      mcause <= _GEN_9;
    end
    if (reset) begin // @[Csr.scala 47:26]
      mcycle <= 64'h0; // @[Csr.scala 47:26]
    end else if (csr_rw) begin // @[Csr.scala 118:13]
      if (addr == 12'hb00) begin // @[Csr.scala 119:32]
        if (4'h9 == io_sysop) begin // @[Mux.scala 80:57]
          mcycle <= _wdata_T_5;
        end else begin
          mcycle <= _wdata_T_13;
        end
      end else begin
        mcycle <= _mcycle_T_1; // @[Csr.scala 87:10]
      end
    end else begin
      mcycle <= _mcycle_T_1; // @[Csr.scala 87:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mstatus = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mie = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mtvec = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mscratch = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mepc = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mcause = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mcycle = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Clint(
  input         clock,
  input         reset,
  input  [63:0] io_mstatus,
  input  [63:0] io_mie,
  input         io_cmp_ren,
  input         io_cmp_wen,
  input  [63:0] io_cmp_addr,
  input  [63:0] io_cmp_wdata,
  output [63:0] io_cmp_rdata,
  output        io_time_int
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[Clint.scala 26:26]
  reg [63:0] mtimecmp; // @[Clint.scala 27:26]
  wire [63:0] _mtime_T_1 = mtime + 64'h1; // @[Clint.scala 29:18]
  wire [63:0] _io_cmp_rdata_T_1 = io_cmp_addr == 64'h200bff8 ? mtime : mtimecmp; // @[Clint.scala 36:35]
  assign io_cmp_rdata = io_cmp_ren ? _io_cmp_rdata_T_1 : 64'h0; // @[Clint.scala 36:22]
  assign io_time_int = mtime >= mtimecmp & io_mstatus[3] & io_mie[7]; // @[Clint.scala 34:59]
  always @(posedge clock) begin
    if (reset) begin // @[Clint.scala 26:26]
      mtime <= 64'h0; // @[Clint.scala 26:26]
    end else begin
      mtime <= _mtime_T_1; // @[Clint.scala 29:9]
    end
    if (reset) begin // @[Clint.scala 27:26]
      mtimecmp <= 64'h0; // @[Clint.scala 27:26]
    end else if (io_cmp_wen) begin // @[Clint.scala 30:18]
      mtimecmp <= io_cmp_wdata; // @[Clint.scala 31:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core(
  input         clock,
  input         reset,
  output        io_imem_inst_valid,
  input         io_imem_inst_ready,
  output [31:0] io_imem_inst_addr,
  input  [31:0] io_imem_inst_read,
  output        io_dmem_data_valid,
  input         io_dmem_data_ready,
  output        io_dmem_data_req,
  output [31:0] io_dmem_data_addr,
  output [1:0]  io_dmem_data_size,
  output [7:0]  io_dmem_data_strb,
  input  [63:0] io_dmem_data_read,
  output [63:0] io_dmem_data_write,
  output        io_br_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  fetch_clock; // @[Core.scala 13:21]
  wire  fetch_reset; // @[Core.scala 13:21]
  wire  fetch_io_imem_inst_valid; // @[Core.scala 13:21]
  wire  fetch_io_imem_inst_ready; // @[Core.scala 13:21]
  wire [31:0] fetch_io_imem_inst_addr; // @[Core.scala 13:21]
  wire [31:0] fetch_io_imem_inst_read; // @[Core.scala 13:21]
  wire [31:0] fetch_io_fe_pc; // @[Core.scala 13:21]
  wire [31:0] fetch_io_fe_inst; // @[Core.scala 13:21]
  wire  fetch_io_br_valid; // @[Core.scala 13:21]
  wire  fetch_io_br_taken; // @[Core.scala 13:21]
  wire [31:0] fetch_io_br_target; // @[Core.scala 13:21]
  wire  fetch_io_csr_jmp; // @[Core.scala 13:21]
  wire [31:0] fetch_io_newpc; // @[Core.scala 13:21]
  wire  fetch_io_instr_valid; // @[Core.scala 13:21]
  wire  fetch_io_flush; // @[Core.scala 13:21]
  wire  fetch_io_if_valid_out; // @[Core.scala 13:21]
  wire  fetch_io_if_allow_out; // @[Core.scala 13:21]
  wire  decode_clock; // @[Core.scala 14:22]
  wire  decode_reset; // @[Core.scala 14:22]
  wire [4:0] decode_io_rs1_addr; // @[Core.scala 14:22]
  wire  decode_io_rs1_en; // @[Core.scala 14:22]
  wire [63:0] decode_io_rs1_data; // @[Core.scala 14:22]
  wire [4:0] decode_io_rs2_addr; // @[Core.scala 14:22]
  wire  decode_io_rs2_en; // @[Core.scala 14:22]
  wire [63:0] decode_io_rs2_data; // @[Core.scala 14:22]
  wire [31:0] decode_io_fe_pc; // @[Core.scala 14:22]
  wire [31:0] decode_io_fe_inst; // @[Core.scala 14:22]
  wire [31:0] decode_io_id_pc; // @[Core.scala 14:22]
  wire [31:0] decode_io_id_inst; // @[Core.scala 14:22]
  wire  decode_io_id_wen; // @[Core.scala 14:22]
  wire [4:0] decode_io_id_wdest; // @[Core.scala 14:22]
  wire [63:0] decode_io_id_op1; // @[Core.scala 14:22]
  wire [63:0] decode_io_id_op2; // @[Core.scala 14:22]
  wire [63:0] decode_io_rs2_value; // @[Core.scala 14:22]
  wire  decode_io_mem_stall; // @[Core.scala 14:22]
  wire  decode_io_instr_valid; // @[Core.scala 14:22]
  wire  decode_io_time_int; // @[Core.scala 14:22]
  wire [4:0] decode_io_EX_wdest; // @[Core.scala 14:22]
  wire [4:0] decode_io_WB_wdest; // @[Core.scala 14:22]
  wire [63:0] decode_io_EX_result; // @[Core.scala 14:22]
  wire [63:0] decode_io_WB_result; // @[Core.scala 14:22]
  wire  decode_io_type_w; // @[Core.scala 14:22]
  wire [11:0] decode_io_idop_aluop; // @[Core.scala 14:22]
  wire [6:0] decode_io_idop_loadop; // @[Core.scala 14:22]
  wire [3:0] decode_io_idop_storeop; // @[Core.scala 14:22]
  wire [3:0] decode_io_idop_sysop; // @[Core.scala 14:22]
  wire  decode_io_inst_my; // @[Core.scala 14:22]
  wire  decode_io_skip; // @[Core.scala 14:22]
  wire [63:0] decode_io_print; // @[Core.scala 14:22]
  wire  decode_io_br_valid; // @[Core.scala 14:22]
  wire  decode_io_br_taken; // @[Core.scala 14:22]
  wire [31:0] decode_io_br_target; // @[Core.scala 14:22]
  wire  decode_io_br_stall; // @[Core.scala 14:22]
  wire  decode_io_flush; // @[Core.scala 14:22]
  wire  decode_io_if_allow_out; // @[Core.scala 14:22]
  wire  decode_io_id_valid_out; // @[Core.scala 14:22]
  wire  decode_io_if_valid_out; // @[Core.scala 14:22]
  wire  decode_io_id_allow_out; // @[Core.scala 14:22]
  wire  execution_clock; // @[Core.scala 15:25]
  wire  execution_reset; // @[Core.scala 15:25]
  wire  execution_io_type_w; // @[Core.scala 15:25]
  wire [63:0] execution_io_csr_rdata; // @[Core.scala 15:25]
  wire [11:0] execution_io_idop_aluop; // @[Core.scala 15:25]
  wire [6:0] execution_io_idop_loadop; // @[Core.scala 15:25]
  wire [3:0] execution_io_idop_storeop; // @[Core.scala 15:25]
  wire [3:0] execution_io_idop_sysop; // @[Core.scala 15:25]
  wire [31:0] execution_io_id_pc; // @[Core.scala 15:25]
  wire [31:0] execution_io_id_inst; // @[Core.scala 15:25]
  wire  execution_io_id_wen; // @[Core.scala 15:25]
  wire [4:0] execution_io_id_wdest; // @[Core.scala 15:25]
  wire [63:0] execution_io_id_op1; // @[Core.scala 15:25]
  wire [63:0] execution_io_id_op2; // @[Core.scala 15:25]
  wire [31:0] execution_io_ex_pc; // @[Core.scala 15:25]
  wire [31:0] execution_io_ex_inst; // @[Core.scala 15:25]
  wire  execution_io_ex_wen; // @[Core.scala 15:25]
  wire [4:0] execution_io_ex_wdest; // @[Core.scala 15:25]
  wire [63:0] execution_io_ex_wdata; // @[Core.scala 15:25]
  wire [63:0] execution_io_ex_op1; // @[Core.scala 15:25]
  wire  execution_io_dmem_data_valid; // @[Core.scala 15:25]
  wire  execution_io_dmem_data_ready; // @[Core.scala 15:25]
  wire  execution_io_dmem_data_req; // @[Core.scala 15:25]
  wire [31:0] execution_io_dmem_data_addr; // @[Core.scala 15:25]
  wire [1:0] execution_io_dmem_data_size; // @[Core.scala 15:25]
  wire [7:0] execution_io_dmem_data_strb; // @[Core.scala 15:25]
  wire [63:0] execution_io_dmem_data_read; // @[Core.scala 15:25]
  wire [63:0] execution_io_dmem_data_write; // @[Core.scala 15:25]
  wire [63:0] execution_io_rs2_value; // @[Core.scala 15:25]
  wire [3:0] execution_io_ex_sysop; // @[Core.scala 15:25]
  wire  execution_io_id_skip; // @[Core.scala 15:25]
  wire  execution_io_cmp_ren; // @[Core.scala 15:25]
  wire  execution_io_cmp_wen; // @[Core.scala 15:25]
  wire [63:0] execution_io_cmp_addr; // @[Core.scala 15:25]
  wire [63:0] execution_io_cmp_wdata; // @[Core.scala 15:25]
  wire [63:0] execution_io_cmp_rdata; // @[Core.scala 15:25]
  wire  execution_io_flush; // @[Core.scala 15:25]
  wire  execution_io_skip; // @[Core.scala 15:25]
  wire  execution_io_mem_stall; // @[Core.scala 15:25]
  wire [4:0] execution_io_EX_wdest; // @[Core.scala 15:25]
  wire [63:0] execution_io_EX_result; // @[Core.scala 15:25]
  wire  execution_io_id_allow_out; // @[Core.scala 15:25]
  wire  execution_io_ex_valid_out; // @[Core.scala 15:25]
  wire  execution_io_id_valid_out; // @[Core.scala 15:25]
  wire  execution_io_ex_allow_out; // @[Core.scala 15:25]
  wire  writeback_clock; // @[Core.scala 16:25]
  wire  writeback_reset; // @[Core.scala 16:25]
  wire [31:0] writeback_io_ex_pc; // @[Core.scala 16:25]
  wire [31:0] writeback_io_ex_inst; // @[Core.scala 16:25]
  wire  writeback_io_ex_wen; // @[Core.scala 16:25]
  wire [4:0] writeback_io_ex_wdest; // @[Core.scala 16:25]
  wire [63:0] writeback_io_ex_wdata; // @[Core.scala 16:25]
  wire [63:0] writeback_io_ex_op1; // @[Core.scala 16:25]
  wire [31:0] writeback_io_wb_pc; // @[Core.scala 16:25]
  wire [31:0] writeback_io_wb_inst; // @[Core.scala 16:25]
  wire  writeback_io_wb_wen; // @[Core.scala 16:25]
  wire [4:0] writeback_io_wb_wdest; // @[Core.scala 16:25]
  wire [63:0] writeback_io_wb_wdata; // @[Core.scala 16:25]
  wire [63:0] writeback_io_wb_op1; // @[Core.scala 16:25]
  wire [3:0] writeback_io_ex_sysop; // @[Core.scala 16:25]
  wire [3:0] writeback_io_sysop; // @[Core.scala 16:25]
  wire  writeback_io_ex_skip; // @[Core.scala 16:25]
  wire  writeback_io_skip; // @[Core.scala 16:25]
  wire  writeback_io_flush; // @[Core.scala 16:25]
  wire  writeback_io_ready_cmt; // @[Core.scala 16:25]
  wire [4:0] writeback_io_WB_wdest; // @[Core.scala 16:25]
  wire [63:0] writeback_io_WB_result; // @[Core.scala 16:25]
  wire  writeback_io_intr; // @[Core.scala 16:25]
  wire  writeback_io_ex_allow_out; // @[Core.scala 16:25]
  wire  writeback_io_ex_valid_out; // @[Core.scala 16:25]
  wire  rf_clock; // @[Core.scala 17:18]
  wire  rf_reset; // @[Core.scala 17:18]
  wire [4:0] rf_io_rs1_addr; // @[Core.scala 17:18]
  wire [4:0] rf_io_rs2_addr; // @[Core.scala 17:18]
  wire [63:0] rf_io_rs1_data; // @[Core.scala 17:18]
  wire [63:0] rf_io_rs2_data; // @[Core.scala 17:18]
  wire [4:0] rf_io_rd_addr; // @[Core.scala 17:18]
  wire [63:0] rf_io_rd_data; // @[Core.scala 17:18]
  wire  rf_io_rd_en; // @[Core.scala 17:18]
  wire [63:0] rf_rf_10; // @[Core.scala 17:18]
  wire  csr_clock; // @[Core.scala 18:19]
  wire  csr_reset; // @[Core.scala 18:19]
  wire [63:0] csr_io_in1; // @[Core.scala 18:19]
  wire [31:0] csr_io_pc; // @[Core.scala 18:19]
  wire [31:0] csr_io_inst; // @[Core.scala 18:19]
  wire [3:0] csr_io_sysop; // @[Core.scala 18:19]
  wire [63:0] csr_io_csr_rdata; // @[Core.scala 18:19]
  wire  csr_io_csr_jmp; // @[Core.scala 18:19]
  wire [31:0] csr_io_newpc; // @[Core.scala 18:19]
  wire [63:0] csr_io_mstatus; // @[Core.scala 18:19]
  wire [63:0] csr_io_mie; // @[Core.scala 18:19]
  wire  csr_io_flush; // @[Core.scala 18:19]
  wire  clint_clock; // @[Core.scala 19:21]
  wire  clint_reset; // @[Core.scala 19:21]
  wire [63:0] clint_io_mstatus; // @[Core.scala 19:21]
  wire [63:0] clint_io_mie; // @[Core.scala 19:21]
  wire  clint_io_cmp_ren; // @[Core.scala 19:21]
  wire  clint_io_cmp_wen; // @[Core.scala 19:21]
  wire [63:0] clint_io_cmp_addr; // @[Core.scala 19:21]
  wire [63:0] clint_io_cmp_wdata; // @[Core.scala 19:21]
  wire [63:0] clint_io_cmp_rdata; // @[Core.scala 19:21]
  wire  clint_io_time_int; // @[Core.scala 19:21]
  wire  dt_ic_clock; // @[Core.scala 108:23]
  wire [7:0] dt_ic_coreid; // @[Core.scala 108:23]
  wire [7:0] dt_ic_index; // @[Core.scala 108:23]
  wire  dt_ic_valid; // @[Core.scala 108:23]
  wire [63:0] dt_ic_pc; // @[Core.scala 108:23]
  wire [31:0] dt_ic_instr; // @[Core.scala 108:23]
  wire [7:0] dt_ic_special; // @[Core.scala 108:23]
  wire  dt_ic_skip; // @[Core.scala 108:23]
  wire  dt_ic_isRVC; // @[Core.scala 108:23]
  wire  dt_ic_scFailed; // @[Core.scala 108:23]
  wire  dt_ic_wen; // @[Core.scala 108:23]
  wire [63:0] dt_ic_wdata; // @[Core.scala 108:23]
  wire [7:0] dt_ic_wdest; // @[Core.scala 108:23]
  wire  dt_ae_clock; // @[Core.scala 123:23]
  wire [7:0] dt_ae_coreid; // @[Core.scala 123:23]
  wire [31:0] dt_ae_intrNO; // @[Core.scala 123:23]
  wire [31:0] dt_ae_cause; // @[Core.scala 123:23]
  wire [63:0] dt_ae_exceptionPC; // @[Core.scala 123:23]
  wire [31:0] dt_ae_exceptionInst; // @[Core.scala 123:23]
  wire  dt_te_clock; // @[Core.scala 139:23]
  wire [7:0] dt_te_coreid; // @[Core.scala 139:23]
  wire  dt_te_valid; // @[Core.scala 139:23]
  wire [2:0] dt_te_code; // @[Core.scala 139:23]
  wire [63:0] dt_te_pc; // @[Core.scala 139:23]
  wire [63:0] dt_te_cycleCnt; // @[Core.scala 139:23]
  wire [63:0] dt_te_instrCnt; // @[Core.scala 139:23]
  reg  inst_my; // @[Core.scala 21:24]
  reg [63:0] print; // @[Core.scala 22:24]
  reg  dt_ic_io_valid_REG; // @[Core.scala 112:33]
  reg [31:0] dt_ic_io_pc_REG; // @[Core.scala 113:33]
  reg [31:0] dt_ic_io_instr_REG; // @[Core.scala 114:33]
  reg  dt_ic_io_skip_REG; // @[Core.scala 116:33]
  reg  dt_ic_io_wen_REG; // @[Core.scala 119:33]
  reg [63:0] dt_ic_io_wdata_REG; // @[Core.scala 120:33]
  reg [4:0] dt_ic_io_wdest_REG; // @[Core.scala 121:33]
  reg [63:0] dt_ae_io_intrNO_REG; // @[Core.scala 126:37]
  reg [31:0] dt_ae_io_exceptionPC_REG; // @[Core.scala 128:37]
  reg [63:0] cycle_cnt; // @[Core.scala 130:28]
  reg [63:0] instr_cnt; // @[Core.scala 131:28]
  wire [63:0] _cycle_cnt_T_1 = cycle_cnt + 64'h1; // @[Core.scala 133:28]
  wire [63:0] _GEN_1 = {{63'd0}, writeback_io_ready_cmt}; // @[Core.scala 134:28]
  wire [63:0] _instr_cnt_T_1 = instr_cnt + _GEN_1; // @[Core.scala 134:28]
  wire [63:0] rf_a0_0 = rf_rf_10;
  InstFetch fetch ( // @[Core.scala 13:21]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_imem_inst_valid(fetch_io_imem_inst_valid),
    .io_imem_inst_ready(fetch_io_imem_inst_ready),
    .io_imem_inst_addr(fetch_io_imem_inst_addr),
    .io_imem_inst_read(fetch_io_imem_inst_read),
    .io_fe_pc(fetch_io_fe_pc),
    .io_fe_inst(fetch_io_fe_inst),
    .io_br_valid(fetch_io_br_valid),
    .io_br_taken(fetch_io_br_taken),
    .io_br_target(fetch_io_br_target),
    .io_csr_jmp(fetch_io_csr_jmp),
    .io_newpc(fetch_io_newpc),
    .io_instr_valid(fetch_io_instr_valid),
    .io_flush(fetch_io_flush),
    .io_if_valid_out(fetch_io_if_valid_out),
    .io_if_allow_out(fetch_io_if_allow_out)
  );
  Decode decode ( // @[Core.scala 14:22]
    .clock(decode_clock),
    .reset(decode_reset),
    .io_rs1_addr(decode_io_rs1_addr),
    .io_rs1_en(decode_io_rs1_en),
    .io_rs1_data(decode_io_rs1_data),
    .io_rs2_addr(decode_io_rs2_addr),
    .io_rs2_en(decode_io_rs2_en),
    .io_rs2_data(decode_io_rs2_data),
    .io_fe_pc(decode_io_fe_pc),
    .io_fe_inst(decode_io_fe_inst),
    .io_id_pc(decode_io_id_pc),
    .io_id_inst(decode_io_id_inst),
    .io_id_wen(decode_io_id_wen),
    .io_id_wdest(decode_io_id_wdest),
    .io_id_op1(decode_io_id_op1),
    .io_id_op2(decode_io_id_op2),
    .io_rs2_value(decode_io_rs2_value),
    .io_mem_stall(decode_io_mem_stall),
    .io_instr_valid(decode_io_instr_valid),
    .io_time_int(decode_io_time_int),
    .io_EX_wdest(decode_io_EX_wdest),
    .io_WB_wdest(decode_io_WB_wdest),
    .io_EX_result(decode_io_EX_result),
    .io_WB_result(decode_io_WB_result),
    .io_type_w(decode_io_type_w),
    .io_idop_aluop(decode_io_idop_aluop),
    .io_idop_loadop(decode_io_idop_loadop),
    .io_idop_storeop(decode_io_idop_storeop),
    .io_idop_sysop(decode_io_idop_sysop),
    .io_inst_my(decode_io_inst_my),
    .io_skip(decode_io_skip),
    .io_print(decode_io_print),
    .io_br_valid(decode_io_br_valid),
    .io_br_taken(decode_io_br_taken),
    .io_br_target(decode_io_br_target),
    .io_br_stall(decode_io_br_stall),
    .io_flush(decode_io_flush),
    .io_if_allow_out(decode_io_if_allow_out),
    .io_id_valid_out(decode_io_id_valid_out),
    .io_if_valid_out(decode_io_if_valid_out),
    .io_id_allow_out(decode_io_id_allow_out)
  );
  Execution execution ( // @[Core.scala 15:25]
    .clock(execution_clock),
    .reset(execution_reset),
    .io_type_w(execution_io_type_w),
    .io_csr_rdata(execution_io_csr_rdata),
    .io_idop_aluop(execution_io_idop_aluop),
    .io_idop_loadop(execution_io_idop_loadop),
    .io_idop_storeop(execution_io_idop_storeop),
    .io_idop_sysop(execution_io_idop_sysop),
    .io_id_pc(execution_io_id_pc),
    .io_id_inst(execution_io_id_inst),
    .io_id_wen(execution_io_id_wen),
    .io_id_wdest(execution_io_id_wdest),
    .io_id_op1(execution_io_id_op1),
    .io_id_op2(execution_io_id_op2),
    .io_ex_pc(execution_io_ex_pc),
    .io_ex_inst(execution_io_ex_inst),
    .io_ex_wen(execution_io_ex_wen),
    .io_ex_wdest(execution_io_ex_wdest),
    .io_ex_wdata(execution_io_ex_wdata),
    .io_ex_op1(execution_io_ex_op1),
    .io_dmem_data_valid(execution_io_dmem_data_valid),
    .io_dmem_data_ready(execution_io_dmem_data_ready),
    .io_dmem_data_req(execution_io_dmem_data_req),
    .io_dmem_data_addr(execution_io_dmem_data_addr),
    .io_dmem_data_size(execution_io_dmem_data_size),
    .io_dmem_data_strb(execution_io_dmem_data_strb),
    .io_dmem_data_read(execution_io_dmem_data_read),
    .io_dmem_data_write(execution_io_dmem_data_write),
    .io_rs2_value(execution_io_rs2_value),
    .io_ex_sysop(execution_io_ex_sysop),
    .io_id_skip(execution_io_id_skip),
    .io_cmp_ren(execution_io_cmp_ren),
    .io_cmp_wen(execution_io_cmp_wen),
    .io_cmp_addr(execution_io_cmp_addr),
    .io_cmp_wdata(execution_io_cmp_wdata),
    .io_cmp_rdata(execution_io_cmp_rdata),
    .io_flush(execution_io_flush),
    .io_skip(execution_io_skip),
    .io_mem_stall(execution_io_mem_stall),
    .io_EX_wdest(execution_io_EX_wdest),
    .io_EX_result(execution_io_EX_result),
    .io_id_allow_out(execution_io_id_allow_out),
    .io_ex_valid_out(execution_io_ex_valid_out),
    .io_id_valid_out(execution_io_id_valid_out),
    .io_ex_allow_out(execution_io_ex_allow_out)
  );
  WriteBack writeback ( // @[Core.scala 16:25]
    .clock(writeback_clock),
    .reset(writeback_reset),
    .io_ex_pc(writeback_io_ex_pc),
    .io_ex_inst(writeback_io_ex_inst),
    .io_ex_wen(writeback_io_ex_wen),
    .io_ex_wdest(writeback_io_ex_wdest),
    .io_ex_wdata(writeback_io_ex_wdata),
    .io_ex_op1(writeback_io_ex_op1),
    .io_wb_pc(writeback_io_wb_pc),
    .io_wb_inst(writeback_io_wb_inst),
    .io_wb_wen(writeback_io_wb_wen),
    .io_wb_wdest(writeback_io_wb_wdest),
    .io_wb_wdata(writeback_io_wb_wdata),
    .io_wb_op1(writeback_io_wb_op1),
    .io_ex_sysop(writeback_io_ex_sysop),
    .io_sysop(writeback_io_sysop),
    .io_ex_skip(writeback_io_ex_skip),
    .io_skip(writeback_io_skip),
    .io_flush(writeback_io_flush),
    .io_ready_cmt(writeback_io_ready_cmt),
    .io_WB_wdest(writeback_io_WB_wdest),
    .io_WB_result(writeback_io_WB_result),
    .io_intr(writeback_io_intr),
    .io_ex_allow_out(writeback_io_ex_allow_out),
    .io_ex_valid_out(writeback_io_ex_valid_out)
  );
  RegFile rf ( // @[Core.scala 17:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_rs1_addr(rf_io_rs1_addr),
    .io_rs2_addr(rf_io_rs2_addr),
    .io_rs1_data(rf_io_rs1_data),
    .io_rs2_data(rf_io_rs2_data),
    .io_rd_addr(rf_io_rd_addr),
    .io_rd_data(rf_io_rd_data),
    .io_rd_en(rf_io_rd_en),
    .rf_10(rf_rf_10)
  );
  Csr csr ( // @[Core.scala 18:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in1(csr_io_in1),
    .io_pc(csr_io_pc),
    .io_inst(csr_io_inst),
    .io_sysop(csr_io_sysop),
    .io_csr_rdata(csr_io_csr_rdata),
    .io_csr_jmp(csr_io_csr_jmp),
    .io_newpc(csr_io_newpc),
    .io_mstatus(csr_io_mstatus),
    .io_mie(csr_io_mie),
    .io_flush(csr_io_flush)
  );
  Clint clint ( // @[Core.scala 19:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io_mstatus(clint_io_mstatus),
    .io_mie(clint_io_mie),
    .io_cmp_ren(clint_io_cmp_ren),
    .io_cmp_wen(clint_io_cmp_wen),
    .io_cmp_addr(clint_io_cmp_addr),
    .io_cmp_wdata(clint_io_cmp_wdata),
    .io_cmp_rdata(clint_io_cmp_rdata),
    .io_time_int(clint_io_time_int)
  );
  DifftestInstrCommit dt_ic ( // @[Core.scala 108:23]
    .clock(dt_ic_clock),
    .coreid(dt_ic_coreid),
    .index(dt_ic_index),
    .valid(dt_ic_valid),
    .pc(dt_ic_pc),
    .instr(dt_ic_instr),
    .special(dt_ic_special),
    .skip(dt_ic_skip),
    .isRVC(dt_ic_isRVC),
    .scFailed(dt_ic_scFailed),
    .wen(dt_ic_wen),
    .wdata(dt_ic_wdata),
    .wdest(dt_ic_wdest)
  );
  DifftestArchEvent dt_ae ( // @[Core.scala 123:23]
    .clock(dt_ae_clock),
    .coreid(dt_ae_coreid),
    .intrNO(dt_ae_intrNO),
    .cause(dt_ae_cause),
    .exceptionPC(dt_ae_exceptionPC),
    .exceptionInst(dt_ae_exceptionInst)
  );
  DifftestTrapEvent dt_te ( // @[Core.scala 139:23]
    .clock(dt_te_clock),
    .coreid(dt_te_coreid),
    .valid(dt_te_valid),
    .code(dt_te_code),
    .pc(dt_te_pc),
    .cycleCnt(dt_te_cycleCnt),
    .instrCnt(dt_te_instrCnt)
  );
  assign io_imem_inst_valid = fetch_io_imem_inst_valid; // @[Core.scala 28:29]
  assign io_imem_inst_addr = fetch_io_imem_inst_addr; // @[Core.scala 28:29]
  assign io_dmem_data_valid = execution_io_dmem_data_valid; // @[Core.scala 54:29]
  assign io_dmem_data_req = execution_io_dmem_data_req; // @[Core.scala 54:29]
  assign io_dmem_data_addr = execution_io_dmem_data_addr; // @[Core.scala 54:29]
  assign io_dmem_data_size = execution_io_dmem_data_size; // @[Core.scala 54:29]
  assign io_dmem_data_strb = execution_io_dmem_data_strb; // @[Core.scala 54:29]
  assign io_dmem_data_write = execution_io_dmem_data_write; // @[Core.scala 54:29]
  assign io_br_stall = decode_io_br_stall; // @[Core.scala 25:15]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_imem_inst_ready = io_imem_inst_ready; // @[Core.scala 28:29]
  assign fetch_io_imem_inst_read = io_imem_inst_read; // @[Core.scala 28:29]
  assign fetch_io_br_valid = decode_io_br_valid; // @[Core.scala 29:29]
  assign fetch_io_br_taken = decode_io_br_taken; // @[Core.scala 30:29]
  assign fetch_io_br_target = decode_io_br_target; // @[Core.scala 31:29]
  assign fetch_io_csr_jmp = csr_io_csr_jmp; // @[Core.scala 32:29]
  assign fetch_io_newpc = csr_io_newpc; // @[Core.scala 33:29]
  assign fetch_io_flush = writeback_io_flush; // @[Core.scala 34:29]
  assign fetch_io_if_allow_out = decode_io_if_allow_out; // @[Core.scala 35:29]
  assign decode_clock = clock;
  assign decode_reset = reset;
  assign decode_io_rs1_data = rf_io_rs1_data; // @[Core.scala 38:29]
  assign decode_io_rs2_data = rf_io_rs2_data; // @[Core.scala 39:29]
  assign decode_io_fe_pc = fetch_io_fe_pc; // @[Core.scala 42:29]
  assign decode_io_fe_inst = fetch_io_fe_inst; // @[Core.scala 42:29]
  assign decode_io_mem_stall = execution_io_mem_stall; // @[Core.scala 43:29]
  assign decode_io_instr_valid = fetch_io_instr_valid; // @[Core.scala 44:29]
  assign decode_io_time_int = clint_io_time_int; // @[Core.scala 52:29]
  assign decode_io_EX_wdest = execution_io_EX_wdest; // @[Core.scala 45:29]
  assign decode_io_WB_wdest = writeback_io_WB_wdest; // @[Core.scala 47:29]
  assign decode_io_EX_result = execution_io_EX_result; // @[Core.scala 46:29]
  assign decode_io_WB_result = writeback_io_WB_result; // @[Core.scala 48:29]
  assign decode_io_flush = writeback_io_flush; // @[Core.scala 49:29]
  assign decode_io_if_valid_out = fetch_io_if_valid_out; // @[Core.scala 40:29]
  assign decode_io_id_allow_out = execution_io_id_allow_out; // @[Core.scala 41:29]
  assign execution_clock = clock;
  assign execution_reset = reset;
  assign execution_io_type_w = decode_io_type_w; // @[Core.scala 55:29]
  assign execution_io_csr_rdata = csr_io_csr_rdata; // @[Core.scala 56:29]
  assign execution_io_idop_aluop = decode_io_idop_aluop; // @[Core.scala 58:29]
  assign execution_io_idop_loadop = decode_io_idop_loadop; // @[Core.scala 58:29]
  assign execution_io_idop_storeop = decode_io_idop_storeop; // @[Core.scala 58:29]
  assign execution_io_idop_sysop = decode_io_idop_sysop; // @[Core.scala 58:29]
  assign execution_io_id_pc = decode_io_id_pc; // @[Core.scala 59:29]
  assign execution_io_id_inst = decode_io_id_inst; // @[Core.scala 59:29]
  assign execution_io_id_wen = decode_io_id_wen; // @[Core.scala 59:29]
  assign execution_io_id_wdest = decode_io_id_wdest; // @[Core.scala 59:29]
  assign execution_io_id_op1 = decode_io_id_op1; // @[Core.scala 59:29]
  assign execution_io_id_op2 = decode_io_id_op2; // @[Core.scala 59:29]
  assign execution_io_dmem_data_ready = io_dmem_data_ready; // @[Core.scala 54:29]
  assign execution_io_dmem_data_read = io_dmem_data_read; // @[Core.scala 54:29]
  assign execution_io_rs2_value = decode_io_rs2_value; // @[Core.scala 60:29]
  assign execution_io_id_skip = decode_io_skip; // @[Core.scala 63:29]
  assign execution_io_cmp_rdata = clint_io_cmp_rdata; // @[Core.scala 57:29]
  assign execution_io_flush = writeback_io_flush; // @[Core.scala 64:29]
  assign execution_io_id_valid_out = decode_io_id_valid_out; // @[Core.scala 61:29]
  assign execution_io_ex_allow_out = writeback_io_ex_allow_out; // @[Core.scala 62:29]
  assign writeback_clock = clock;
  assign writeback_reset = reset;
  assign writeback_io_ex_pc = execution_io_ex_pc; // @[Core.scala 67:29]
  assign writeback_io_ex_inst = execution_io_ex_inst; // @[Core.scala 67:29]
  assign writeback_io_ex_wen = execution_io_ex_wen; // @[Core.scala 67:29]
  assign writeback_io_ex_wdest = execution_io_ex_wdest; // @[Core.scala 67:29]
  assign writeback_io_ex_wdata = execution_io_ex_wdata; // @[Core.scala 67:29]
  assign writeback_io_ex_op1 = execution_io_ex_op1; // @[Core.scala 67:29]
  assign writeback_io_ex_sysop = execution_io_ex_sysop; // @[Core.scala 66:29]
  assign writeback_io_ex_skip = execution_io_skip; // @[Core.scala 69:29]
  assign writeback_io_ex_valid_out = execution_io_ex_valid_out; // @[Core.scala 68:29]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_rs1_addr = decode_io_rs1_addr; // @[Core.scala 71:29]
  assign rf_io_rs2_addr = decode_io_rs2_addr; // @[Core.scala 72:29]
  assign rf_io_rd_addr = writeback_io_wb_wdest; // @[Core.scala 73:29]
  assign rf_io_rd_data = writeback_io_wb_wdata; // @[Core.scala 75:29]
  assign rf_io_rd_en = writeback_io_wb_wen; // @[Core.scala 74:29]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in1 = writeback_io_wb_op1; // @[Core.scala 77:29]
  assign csr_io_pc = writeback_io_wb_pc; // @[Core.scala 80:29]
  assign csr_io_inst = execution_io_ex_inst; // @[Core.scala 79:29]
  assign csr_io_sysop = writeback_io_sysop; // @[Core.scala 78:29]
  assign csr_io_flush = writeback_io_flush; // @[Core.scala 81:29]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io_mstatus = csr_io_mstatus; // @[Core.scala 83:29]
  assign clint_io_mie = csr_io_mie; // @[Core.scala 84:29]
  assign clint_io_cmp_ren = execution_io_cmp_ren; // @[Core.scala 85:29]
  assign clint_io_cmp_wen = execution_io_cmp_wen; // @[Core.scala 86:29]
  assign clint_io_cmp_addr = execution_io_cmp_addr; // @[Core.scala 87:29]
  assign clint_io_cmp_wdata = execution_io_cmp_wdata; // @[Core.scala 88:29]
  assign dt_ic_clock = clock; // @[Core.scala 109:23]
  assign dt_ic_coreid = 8'h0; // @[Core.scala 110:23]
  assign dt_ic_index = 8'h0; // @[Core.scala 111:23]
  assign dt_ic_valid = dt_ic_io_valid_REG; // @[Core.scala 112:23]
  assign dt_ic_pc = {{32'd0}, dt_ic_io_pc_REG}; // @[Core.scala 113:23]
  assign dt_ic_instr = dt_ic_io_instr_REG; // @[Core.scala 114:23]
  assign dt_ic_special = 8'h0; // @[Core.scala 115:23]
  assign dt_ic_skip = dt_ic_io_skip_REG; // @[Core.scala 116:23]
  assign dt_ic_isRVC = 1'h0; // @[Core.scala 117:23]
  assign dt_ic_scFailed = 1'h0; // @[Core.scala 118:23]
  assign dt_ic_wen = dt_ic_io_wen_REG; // @[Core.scala 119:23]
  assign dt_ic_wdata = dt_ic_io_wdata_REG; // @[Core.scala 120:23]
  assign dt_ic_wdest = {{3'd0}, dt_ic_io_wdest_REG}; // @[Core.scala 121:23]
  assign dt_ae_clock = clock; // @[Core.scala 124:27]
  assign dt_ae_coreid = 8'h0; // @[Core.scala 125:27]
  assign dt_ae_intrNO = dt_ae_io_intrNO_REG[31:0]; // @[Core.scala 126:27]
  assign dt_ae_cause = 32'h0; // @[Core.scala 127:27]
  assign dt_ae_exceptionPC = {{32'd0}, dt_ae_io_exceptionPC_REG}; // @[Core.scala 128:27]
  assign dt_ae_exceptionInst = 32'h0;
  assign dt_te_clock = clock; // @[Core.scala 140:23]
  assign dt_te_coreid = 8'h0; // @[Core.scala 141:23]
  assign dt_te_valid = writeback_io_wb_inst == 32'h6b; // @[Core.scala 142:48]
  assign dt_te_code = rf_a0_0[2:0]; // @[Core.scala 143:31]
  assign dt_te_pc = {{32'd0}, writeback_io_wb_pc}; // @[Core.scala 144:23]
  assign dt_te_cycleCnt = cycle_cnt; // @[Core.scala 145:23]
  assign dt_te_instrCnt = instr_cnt; // @[Core.scala 146:23]
  always @(posedge clock) begin
    if (reset) begin // @[Core.scala 21:24]
      inst_my <= 1'h0; // @[Core.scala 21:24]
    end else begin
      inst_my <= decode_io_inst_my; // @[Core.scala 95:11]
    end
    if (reset) begin // @[Core.scala 22:24]
      print <= 64'h0; // @[Core.scala 22:24]
    end else if (inst_my) begin // @[Core.scala 96:18]
      print <= decode_io_print; // @[Core.scala 97:11]
    end
    dt_ic_io_valid_REG <= writeback_io_ready_cmt; // @[Core.scala 112:33]
    dt_ic_io_pc_REG <= writeback_io_wb_pc; // @[Core.scala 113:33]
    dt_ic_io_instr_REG <= writeback_io_wb_inst; // @[Core.scala 114:33]
    dt_ic_io_skip_REG <= writeback_io_skip | csr_io_inst[31:20] == 12'hb00 & csr_io_sysop != 4'h0; // @[Core.scala 23:35]
    dt_ic_io_wen_REG <= writeback_io_wb_wen; // @[Core.scala 119:33]
    dt_ic_io_wdata_REG <= writeback_io_wb_wdata; // @[Core.scala 120:33]
    dt_ic_io_wdest_REG <= writeback_io_wb_wdest; // @[Core.scala 121:33]
    if (writeback_io_intr) begin // @[Core.scala 104:20]
      dt_ae_io_intrNO_REG <= 64'h7;
    end else begin
      dt_ae_io_intrNO_REG <= 64'h0;
    end
    if (writeback_io_intr) begin // @[Core.scala 105:24]
      dt_ae_io_exceptionPC_REG <= writeback_io_wb_pc;
    end else begin
      dt_ae_io_exceptionPC_REG <= 32'h0;
    end
    if (reset) begin // @[Core.scala 130:28]
      cycle_cnt <= 64'h0; // @[Core.scala 130:28]
    end else begin
      cycle_cnt <= _cycle_cnt_T_1; // @[Core.scala 133:15]
    end
    if (reset) begin // @[Core.scala 131:28]
      instr_cnt <= 64'h0; // @[Core.scala 131:28]
    end else begin
      instr_cnt <= _instr_cnt_T_1; // @[Core.scala 134:15]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (writeback_io_ready_cmt & ~reset) begin
          $fwrite(32'h80000002,"%c",print); // @[Core.scala 100:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst_my = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  print = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  dt_ic_io_valid_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  dt_ic_io_pc_REG = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  dt_ic_io_instr_REG = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  dt_ic_io_skip_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dt_ic_io_wen_REG = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  dt_ic_io_wdata_REG = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  dt_ic_io_wdest_REG = _RAND_8[4:0];
  _RAND_9 = {2{`RANDOM}};
  dt_ae_io_intrNO_REG = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  dt_ae_io_exceptionPC_REG = _RAND_10[31:0];
  _RAND_11 = {2{`RANDOM}};
  cycle_cnt = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  instr_cnt = _RAND_12[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Icache(
  input          clock,
  input          reset,
  input          io_imem_inst_valid,
  output         io_imem_inst_ready,
  input  [31:0]  io_imem_inst_addr,
  output [31:0]  io_imem_inst_read,
  output         io_out_inst_valid,
  input          io_out_inst_ready,
  output [31:0]  io_out_inst_addr,
  input  [127:0] io_out_inst_read,
  input          io_br_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [127:0] _RAND_516;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] req_Q; // @[Icache.scala 126:19]
  wire  req_CLK; // @[Icache.scala 126:19]
  wire  req_CEN; // @[Icache.scala 126:19]
  wire  req_WEN; // @[Icache.scala 126:19]
  wire [7:0] req_A; // @[Icache.scala 126:19]
  wire [127:0] req_D; // @[Icache.scala 126:19]
  reg [19:0] tag_0; // @[Icache.scala 17:24]
  reg [19:0] tag_1; // @[Icache.scala 17:24]
  reg [19:0] tag_2; // @[Icache.scala 17:24]
  reg [19:0] tag_3; // @[Icache.scala 17:24]
  reg [19:0] tag_4; // @[Icache.scala 17:24]
  reg [19:0] tag_5; // @[Icache.scala 17:24]
  reg [19:0] tag_6; // @[Icache.scala 17:24]
  reg [19:0] tag_7; // @[Icache.scala 17:24]
  reg [19:0] tag_8; // @[Icache.scala 17:24]
  reg [19:0] tag_9; // @[Icache.scala 17:24]
  reg [19:0] tag_10; // @[Icache.scala 17:24]
  reg [19:0] tag_11; // @[Icache.scala 17:24]
  reg [19:0] tag_12; // @[Icache.scala 17:24]
  reg [19:0] tag_13; // @[Icache.scala 17:24]
  reg [19:0] tag_14; // @[Icache.scala 17:24]
  reg [19:0] tag_15; // @[Icache.scala 17:24]
  reg [19:0] tag_16; // @[Icache.scala 17:24]
  reg [19:0] tag_17; // @[Icache.scala 17:24]
  reg [19:0] tag_18; // @[Icache.scala 17:24]
  reg [19:0] tag_19; // @[Icache.scala 17:24]
  reg [19:0] tag_20; // @[Icache.scala 17:24]
  reg [19:0] tag_21; // @[Icache.scala 17:24]
  reg [19:0] tag_22; // @[Icache.scala 17:24]
  reg [19:0] tag_23; // @[Icache.scala 17:24]
  reg [19:0] tag_24; // @[Icache.scala 17:24]
  reg [19:0] tag_25; // @[Icache.scala 17:24]
  reg [19:0] tag_26; // @[Icache.scala 17:24]
  reg [19:0] tag_27; // @[Icache.scala 17:24]
  reg [19:0] tag_28; // @[Icache.scala 17:24]
  reg [19:0] tag_29; // @[Icache.scala 17:24]
  reg [19:0] tag_30; // @[Icache.scala 17:24]
  reg [19:0] tag_31; // @[Icache.scala 17:24]
  reg [19:0] tag_32; // @[Icache.scala 17:24]
  reg [19:0] tag_33; // @[Icache.scala 17:24]
  reg [19:0] tag_34; // @[Icache.scala 17:24]
  reg [19:0] tag_35; // @[Icache.scala 17:24]
  reg [19:0] tag_36; // @[Icache.scala 17:24]
  reg [19:0] tag_37; // @[Icache.scala 17:24]
  reg [19:0] tag_38; // @[Icache.scala 17:24]
  reg [19:0] tag_39; // @[Icache.scala 17:24]
  reg [19:0] tag_40; // @[Icache.scala 17:24]
  reg [19:0] tag_41; // @[Icache.scala 17:24]
  reg [19:0] tag_42; // @[Icache.scala 17:24]
  reg [19:0] tag_43; // @[Icache.scala 17:24]
  reg [19:0] tag_44; // @[Icache.scala 17:24]
  reg [19:0] tag_45; // @[Icache.scala 17:24]
  reg [19:0] tag_46; // @[Icache.scala 17:24]
  reg [19:0] tag_47; // @[Icache.scala 17:24]
  reg [19:0] tag_48; // @[Icache.scala 17:24]
  reg [19:0] tag_49; // @[Icache.scala 17:24]
  reg [19:0] tag_50; // @[Icache.scala 17:24]
  reg [19:0] tag_51; // @[Icache.scala 17:24]
  reg [19:0] tag_52; // @[Icache.scala 17:24]
  reg [19:0] tag_53; // @[Icache.scala 17:24]
  reg [19:0] tag_54; // @[Icache.scala 17:24]
  reg [19:0] tag_55; // @[Icache.scala 17:24]
  reg [19:0] tag_56; // @[Icache.scala 17:24]
  reg [19:0] tag_57; // @[Icache.scala 17:24]
  reg [19:0] tag_58; // @[Icache.scala 17:24]
  reg [19:0] tag_59; // @[Icache.scala 17:24]
  reg [19:0] tag_60; // @[Icache.scala 17:24]
  reg [19:0] tag_61; // @[Icache.scala 17:24]
  reg [19:0] tag_62; // @[Icache.scala 17:24]
  reg [19:0] tag_63; // @[Icache.scala 17:24]
  reg [19:0] tag_64; // @[Icache.scala 17:24]
  reg [19:0] tag_65; // @[Icache.scala 17:24]
  reg [19:0] tag_66; // @[Icache.scala 17:24]
  reg [19:0] tag_67; // @[Icache.scala 17:24]
  reg [19:0] tag_68; // @[Icache.scala 17:24]
  reg [19:0] tag_69; // @[Icache.scala 17:24]
  reg [19:0] tag_70; // @[Icache.scala 17:24]
  reg [19:0] tag_71; // @[Icache.scala 17:24]
  reg [19:0] tag_72; // @[Icache.scala 17:24]
  reg [19:0] tag_73; // @[Icache.scala 17:24]
  reg [19:0] tag_74; // @[Icache.scala 17:24]
  reg [19:0] tag_75; // @[Icache.scala 17:24]
  reg [19:0] tag_76; // @[Icache.scala 17:24]
  reg [19:0] tag_77; // @[Icache.scala 17:24]
  reg [19:0] tag_78; // @[Icache.scala 17:24]
  reg [19:0] tag_79; // @[Icache.scala 17:24]
  reg [19:0] tag_80; // @[Icache.scala 17:24]
  reg [19:0] tag_81; // @[Icache.scala 17:24]
  reg [19:0] tag_82; // @[Icache.scala 17:24]
  reg [19:0] tag_83; // @[Icache.scala 17:24]
  reg [19:0] tag_84; // @[Icache.scala 17:24]
  reg [19:0] tag_85; // @[Icache.scala 17:24]
  reg [19:0] tag_86; // @[Icache.scala 17:24]
  reg [19:0] tag_87; // @[Icache.scala 17:24]
  reg [19:0] tag_88; // @[Icache.scala 17:24]
  reg [19:0] tag_89; // @[Icache.scala 17:24]
  reg [19:0] tag_90; // @[Icache.scala 17:24]
  reg [19:0] tag_91; // @[Icache.scala 17:24]
  reg [19:0] tag_92; // @[Icache.scala 17:24]
  reg [19:0] tag_93; // @[Icache.scala 17:24]
  reg [19:0] tag_94; // @[Icache.scala 17:24]
  reg [19:0] tag_95; // @[Icache.scala 17:24]
  reg [19:0] tag_96; // @[Icache.scala 17:24]
  reg [19:0] tag_97; // @[Icache.scala 17:24]
  reg [19:0] tag_98; // @[Icache.scala 17:24]
  reg [19:0] tag_99; // @[Icache.scala 17:24]
  reg [19:0] tag_100; // @[Icache.scala 17:24]
  reg [19:0] tag_101; // @[Icache.scala 17:24]
  reg [19:0] tag_102; // @[Icache.scala 17:24]
  reg [19:0] tag_103; // @[Icache.scala 17:24]
  reg [19:0] tag_104; // @[Icache.scala 17:24]
  reg [19:0] tag_105; // @[Icache.scala 17:24]
  reg [19:0] tag_106; // @[Icache.scala 17:24]
  reg [19:0] tag_107; // @[Icache.scala 17:24]
  reg [19:0] tag_108; // @[Icache.scala 17:24]
  reg [19:0] tag_109; // @[Icache.scala 17:24]
  reg [19:0] tag_110; // @[Icache.scala 17:24]
  reg [19:0] tag_111; // @[Icache.scala 17:24]
  reg [19:0] tag_112; // @[Icache.scala 17:24]
  reg [19:0] tag_113; // @[Icache.scala 17:24]
  reg [19:0] tag_114; // @[Icache.scala 17:24]
  reg [19:0] tag_115; // @[Icache.scala 17:24]
  reg [19:0] tag_116; // @[Icache.scala 17:24]
  reg [19:0] tag_117; // @[Icache.scala 17:24]
  reg [19:0] tag_118; // @[Icache.scala 17:24]
  reg [19:0] tag_119; // @[Icache.scala 17:24]
  reg [19:0] tag_120; // @[Icache.scala 17:24]
  reg [19:0] tag_121; // @[Icache.scala 17:24]
  reg [19:0] tag_122; // @[Icache.scala 17:24]
  reg [19:0] tag_123; // @[Icache.scala 17:24]
  reg [19:0] tag_124; // @[Icache.scala 17:24]
  reg [19:0] tag_125; // @[Icache.scala 17:24]
  reg [19:0] tag_126; // @[Icache.scala 17:24]
  reg [19:0] tag_127; // @[Icache.scala 17:24]
  reg [19:0] tag_128; // @[Icache.scala 17:24]
  reg [19:0] tag_129; // @[Icache.scala 17:24]
  reg [19:0] tag_130; // @[Icache.scala 17:24]
  reg [19:0] tag_131; // @[Icache.scala 17:24]
  reg [19:0] tag_132; // @[Icache.scala 17:24]
  reg [19:0] tag_133; // @[Icache.scala 17:24]
  reg [19:0] tag_134; // @[Icache.scala 17:24]
  reg [19:0] tag_135; // @[Icache.scala 17:24]
  reg [19:0] tag_136; // @[Icache.scala 17:24]
  reg [19:0] tag_137; // @[Icache.scala 17:24]
  reg [19:0] tag_138; // @[Icache.scala 17:24]
  reg [19:0] tag_139; // @[Icache.scala 17:24]
  reg [19:0] tag_140; // @[Icache.scala 17:24]
  reg [19:0] tag_141; // @[Icache.scala 17:24]
  reg [19:0] tag_142; // @[Icache.scala 17:24]
  reg [19:0] tag_143; // @[Icache.scala 17:24]
  reg [19:0] tag_144; // @[Icache.scala 17:24]
  reg [19:0] tag_145; // @[Icache.scala 17:24]
  reg [19:0] tag_146; // @[Icache.scala 17:24]
  reg [19:0] tag_147; // @[Icache.scala 17:24]
  reg [19:0] tag_148; // @[Icache.scala 17:24]
  reg [19:0] tag_149; // @[Icache.scala 17:24]
  reg [19:0] tag_150; // @[Icache.scala 17:24]
  reg [19:0] tag_151; // @[Icache.scala 17:24]
  reg [19:0] tag_152; // @[Icache.scala 17:24]
  reg [19:0] tag_153; // @[Icache.scala 17:24]
  reg [19:0] tag_154; // @[Icache.scala 17:24]
  reg [19:0] tag_155; // @[Icache.scala 17:24]
  reg [19:0] tag_156; // @[Icache.scala 17:24]
  reg [19:0] tag_157; // @[Icache.scala 17:24]
  reg [19:0] tag_158; // @[Icache.scala 17:24]
  reg [19:0] tag_159; // @[Icache.scala 17:24]
  reg [19:0] tag_160; // @[Icache.scala 17:24]
  reg [19:0] tag_161; // @[Icache.scala 17:24]
  reg [19:0] tag_162; // @[Icache.scala 17:24]
  reg [19:0] tag_163; // @[Icache.scala 17:24]
  reg [19:0] tag_164; // @[Icache.scala 17:24]
  reg [19:0] tag_165; // @[Icache.scala 17:24]
  reg [19:0] tag_166; // @[Icache.scala 17:24]
  reg [19:0] tag_167; // @[Icache.scala 17:24]
  reg [19:0] tag_168; // @[Icache.scala 17:24]
  reg [19:0] tag_169; // @[Icache.scala 17:24]
  reg [19:0] tag_170; // @[Icache.scala 17:24]
  reg [19:0] tag_171; // @[Icache.scala 17:24]
  reg [19:0] tag_172; // @[Icache.scala 17:24]
  reg [19:0] tag_173; // @[Icache.scala 17:24]
  reg [19:0] tag_174; // @[Icache.scala 17:24]
  reg [19:0] tag_175; // @[Icache.scala 17:24]
  reg [19:0] tag_176; // @[Icache.scala 17:24]
  reg [19:0] tag_177; // @[Icache.scala 17:24]
  reg [19:0] tag_178; // @[Icache.scala 17:24]
  reg [19:0] tag_179; // @[Icache.scala 17:24]
  reg [19:0] tag_180; // @[Icache.scala 17:24]
  reg [19:0] tag_181; // @[Icache.scala 17:24]
  reg [19:0] tag_182; // @[Icache.scala 17:24]
  reg [19:0] tag_183; // @[Icache.scala 17:24]
  reg [19:0] tag_184; // @[Icache.scala 17:24]
  reg [19:0] tag_185; // @[Icache.scala 17:24]
  reg [19:0] tag_186; // @[Icache.scala 17:24]
  reg [19:0] tag_187; // @[Icache.scala 17:24]
  reg [19:0] tag_188; // @[Icache.scala 17:24]
  reg [19:0] tag_189; // @[Icache.scala 17:24]
  reg [19:0] tag_190; // @[Icache.scala 17:24]
  reg [19:0] tag_191; // @[Icache.scala 17:24]
  reg [19:0] tag_192; // @[Icache.scala 17:24]
  reg [19:0] tag_193; // @[Icache.scala 17:24]
  reg [19:0] tag_194; // @[Icache.scala 17:24]
  reg [19:0] tag_195; // @[Icache.scala 17:24]
  reg [19:0] tag_196; // @[Icache.scala 17:24]
  reg [19:0] tag_197; // @[Icache.scala 17:24]
  reg [19:0] tag_198; // @[Icache.scala 17:24]
  reg [19:0] tag_199; // @[Icache.scala 17:24]
  reg [19:0] tag_200; // @[Icache.scala 17:24]
  reg [19:0] tag_201; // @[Icache.scala 17:24]
  reg [19:0] tag_202; // @[Icache.scala 17:24]
  reg [19:0] tag_203; // @[Icache.scala 17:24]
  reg [19:0] tag_204; // @[Icache.scala 17:24]
  reg [19:0] tag_205; // @[Icache.scala 17:24]
  reg [19:0] tag_206; // @[Icache.scala 17:24]
  reg [19:0] tag_207; // @[Icache.scala 17:24]
  reg [19:0] tag_208; // @[Icache.scala 17:24]
  reg [19:0] tag_209; // @[Icache.scala 17:24]
  reg [19:0] tag_210; // @[Icache.scala 17:24]
  reg [19:0] tag_211; // @[Icache.scala 17:24]
  reg [19:0] tag_212; // @[Icache.scala 17:24]
  reg [19:0] tag_213; // @[Icache.scala 17:24]
  reg [19:0] tag_214; // @[Icache.scala 17:24]
  reg [19:0] tag_215; // @[Icache.scala 17:24]
  reg [19:0] tag_216; // @[Icache.scala 17:24]
  reg [19:0] tag_217; // @[Icache.scala 17:24]
  reg [19:0] tag_218; // @[Icache.scala 17:24]
  reg [19:0] tag_219; // @[Icache.scala 17:24]
  reg [19:0] tag_220; // @[Icache.scala 17:24]
  reg [19:0] tag_221; // @[Icache.scala 17:24]
  reg [19:0] tag_222; // @[Icache.scala 17:24]
  reg [19:0] tag_223; // @[Icache.scala 17:24]
  reg [19:0] tag_224; // @[Icache.scala 17:24]
  reg [19:0] tag_225; // @[Icache.scala 17:24]
  reg [19:0] tag_226; // @[Icache.scala 17:24]
  reg [19:0] tag_227; // @[Icache.scala 17:24]
  reg [19:0] tag_228; // @[Icache.scala 17:24]
  reg [19:0] tag_229; // @[Icache.scala 17:24]
  reg [19:0] tag_230; // @[Icache.scala 17:24]
  reg [19:0] tag_231; // @[Icache.scala 17:24]
  reg [19:0] tag_232; // @[Icache.scala 17:24]
  reg [19:0] tag_233; // @[Icache.scala 17:24]
  reg [19:0] tag_234; // @[Icache.scala 17:24]
  reg [19:0] tag_235; // @[Icache.scala 17:24]
  reg [19:0] tag_236; // @[Icache.scala 17:24]
  reg [19:0] tag_237; // @[Icache.scala 17:24]
  reg [19:0] tag_238; // @[Icache.scala 17:24]
  reg [19:0] tag_239; // @[Icache.scala 17:24]
  reg [19:0] tag_240; // @[Icache.scala 17:24]
  reg [19:0] tag_241; // @[Icache.scala 17:24]
  reg [19:0] tag_242; // @[Icache.scala 17:24]
  reg [19:0] tag_243; // @[Icache.scala 17:24]
  reg [19:0] tag_244; // @[Icache.scala 17:24]
  reg [19:0] tag_245; // @[Icache.scala 17:24]
  reg [19:0] tag_246; // @[Icache.scala 17:24]
  reg [19:0] tag_247; // @[Icache.scala 17:24]
  reg [19:0] tag_248; // @[Icache.scala 17:24]
  reg [19:0] tag_249; // @[Icache.scala 17:24]
  reg [19:0] tag_250; // @[Icache.scala 17:24]
  reg [19:0] tag_251; // @[Icache.scala 17:24]
  reg [19:0] tag_252; // @[Icache.scala 17:24]
  reg [19:0] tag_253; // @[Icache.scala 17:24]
  reg [19:0] tag_254; // @[Icache.scala 17:24]
  reg [19:0] tag_255; // @[Icache.scala 17:24]
  reg  valid_0; // @[Icache.scala 18:24]
  reg  valid_1; // @[Icache.scala 18:24]
  reg  valid_2; // @[Icache.scala 18:24]
  reg  valid_3; // @[Icache.scala 18:24]
  reg  valid_4; // @[Icache.scala 18:24]
  reg  valid_5; // @[Icache.scala 18:24]
  reg  valid_6; // @[Icache.scala 18:24]
  reg  valid_7; // @[Icache.scala 18:24]
  reg  valid_8; // @[Icache.scala 18:24]
  reg  valid_9; // @[Icache.scala 18:24]
  reg  valid_10; // @[Icache.scala 18:24]
  reg  valid_11; // @[Icache.scala 18:24]
  reg  valid_12; // @[Icache.scala 18:24]
  reg  valid_13; // @[Icache.scala 18:24]
  reg  valid_14; // @[Icache.scala 18:24]
  reg  valid_15; // @[Icache.scala 18:24]
  reg  valid_16; // @[Icache.scala 18:24]
  reg  valid_17; // @[Icache.scala 18:24]
  reg  valid_18; // @[Icache.scala 18:24]
  reg  valid_19; // @[Icache.scala 18:24]
  reg  valid_20; // @[Icache.scala 18:24]
  reg  valid_21; // @[Icache.scala 18:24]
  reg  valid_22; // @[Icache.scala 18:24]
  reg  valid_23; // @[Icache.scala 18:24]
  reg  valid_24; // @[Icache.scala 18:24]
  reg  valid_25; // @[Icache.scala 18:24]
  reg  valid_26; // @[Icache.scala 18:24]
  reg  valid_27; // @[Icache.scala 18:24]
  reg  valid_28; // @[Icache.scala 18:24]
  reg  valid_29; // @[Icache.scala 18:24]
  reg  valid_30; // @[Icache.scala 18:24]
  reg  valid_31; // @[Icache.scala 18:24]
  reg  valid_32; // @[Icache.scala 18:24]
  reg  valid_33; // @[Icache.scala 18:24]
  reg  valid_34; // @[Icache.scala 18:24]
  reg  valid_35; // @[Icache.scala 18:24]
  reg  valid_36; // @[Icache.scala 18:24]
  reg  valid_37; // @[Icache.scala 18:24]
  reg  valid_38; // @[Icache.scala 18:24]
  reg  valid_39; // @[Icache.scala 18:24]
  reg  valid_40; // @[Icache.scala 18:24]
  reg  valid_41; // @[Icache.scala 18:24]
  reg  valid_42; // @[Icache.scala 18:24]
  reg  valid_43; // @[Icache.scala 18:24]
  reg  valid_44; // @[Icache.scala 18:24]
  reg  valid_45; // @[Icache.scala 18:24]
  reg  valid_46; // @[Icache.scala 18:24]
  reg  valid_47; // @[Icache.scala 18:24]
  reg  valid_48; // @[Icache.scala 18:24]
  reg  valid_49; // @[Icache.scala 18:24]
  reg  valid_50; // @[Icache.scala 18:24]
  reg  valid_51; // @[Icache.scala 18:24]
  reg  valid_52; // @[Icache.scala 18:24]
  reg  valid_53; // @[Icache.scala 18:24]
  reg  valid_54; // @[Icache.scala 18:24]
  reg  valid_55; // @[Icache.scala 18:24]
  reg  valid_56; // @[Icache.scala 18:24]
  reg  valid_57; // @[Icache.scala 18:24]
  reg  valid_58; // @[Icache.scala 18:24]
  reg  valid_59; // @[Icache.scala 18:24]
  reg  valid_60; // @[Icache.scala 18:24]
  reg  valid_61; // @[Icache.scala 18:24]
  reg  valid_62; // @[Icache.scala 18:24]
  reg  valid_63; // @[Icache.scala 18:24]
  reg  valid_64; // @[Icache.scala 18:24]
  reg  valid_65; // @[Icache.scala 18:24]
  reg  valid_66; // @[Icache.scala 18:24]
  reg  valid_67; // @[Icache.scala 18:24]
  reg  valid_68; // @[Icache.scala 18:24]
  reg  valid_69; // @[Icache.scala 18:24]
  reg  valid_70; // @[Icache.scala 18:24]
  reg  valid_71; // @[Icache.scala 18:24]
  reg  valid_72; // @[Icache.scala 18:24]
  reg  valid_73; // @[Icache.scala 18:24]
  reg  valid_74; // @[Icache.scala 18:24]
  reg  valid_75; // @[Icache.scala 18:24]
  reg  valid_76; // @[Icache.scala 18:24]
  reg  valid_77; // @[Icache.scala 18:24]
  reg  valid_78; // @[Icache.scala 18:24]
  reg  valid_79; // @[Icache.scala 18:24]
  reg  valid_80; // @[Icache.scala 18:24]
  reg  valid_81; // @[Icache.scala 18:24]
  reg  valid_82; // @[Icache.scala 18:24]
  reg  valid_83; // @[Icache.scala 18:24]
  reg  valid_84; // @[Icache.scala 18:24]
  reg  valid_85; // @[Icache.scala 18:24]
  reg  valid_86; // @[Icache.scala 18:24]
  reg  valid_87; // @[Icache.scala 18:24]
  reg  valid_88; // @[Icache.scala 18:24]
  reg  valid_89; // @[Icache.scala 18:24]
  reg  valid_90; // @[Icache.scala 18:24]
  reg  valid_91; // @[Icache.scala 18:24]
  reg  valid_92; // @[Icache.scala 18:24]
  reg  valid_93; // @[Icache.scala 18:24]
  reg  valid_94; // @[Icache.scala 18:24]
  reg  valid_95; // @[Icache.scala 18:24]
  reg  valid_96; // @[Icache.scala 18:24]
  reg  valid_97; // @[Icache.scala 18:24]
  reg  valid_98; // @[Icache.scala 18:24]
  reg  valid_99; // @[Icache.scala 18:24]
  reg  valid_100; // @[Icache.scala 18:24]
  reg  valid_101; // @[Icache.scala 18:24]
  reg  valid_102; // @[Icache.scala 18:24]
  reg  valid_103; // @[Icache.scala 18:24]
  reg  valid_104; // @[Icache.scala 18:24]
  reg  valid_105; // @[Icache.scala 18:24]
  reg  valid_106; // @[Icache.scala 18:24]
  reg  valid_107; // @[Icache.scala 18:24]
  reg  valid_108; // @[Icache.scala 18:24]
  reg  valid_109; // @[Icache.scala 18:24]
  reg  valid_110; // @[Icache.scala 18:24]
  reg  valid_111; // @[Icache.scala 18:24]
  reg  valid_112; // @[Icache.scala 18:24]
  reg  valid_113; // @[Icache.scala 18:24]
  reg  valid_114; // @[Icache.scala 18:24]
  reg  valid_115; // @[Icache.scala 18:24]
  reg  valid_116; // @[Icache.scala 18:24]
  reg  valid_117; // @[Icache.scala 18:24]
  reg  valid_118; // @[Icache.scala 18:24]
  reg  valid_119; // @[Icache.scala 18:24]
  reg  valid_120; // @[Icache.scala 18:24]
  reg  valid_121; // @[Icache.scala 18:24]
  reg  valid_122; // @[Icache.scala 18:24]
  reg  valid_123; // @[Icache.scala 18:24]
  reg  valid_124; // @[Icache.scala 18:24]
  reg  valid_125; // @[Icache.scala 18:24]
  reg  valid_126; // @[Icache.scala 18:24]
  reg  valid_127; // @[Icache.scala 18:24]
  reg  valid_128; // @[Icache.scala 18:24]
  reg  valid_129; // @[Icache.scala 18:24]
  reg  valid_130; // @[Icache.scala 18:24]
  reg  valid_131; // @[Icache.scala 18:24]
  reg  valid_132; // @[Icache.scala 18:24]
  reg  valid_133; // @[Icache.scala 18:24]
  reg  valid_134; // @[Icache.scala 18:24]
  reg  valid_135; // @[Icache.scala 18:24]
  reg  valid_136; // @[Icache.scala 18:24]
  reg  valid_137; // @[Icache.scala 18:24]
  reg  valid_138; // @[Icache.scala 18:24]
  reg  valid_139; // @[Icache.scala 18:24]
  reg  valid_140; // @[Icache.scala 18:24]
  reg  valid_141; // @[Icache.scala 18:24]
  reg  valid_142; // @[Icache.scala 18:24]
  reg  valid_143; // @[Icache.scala 18:24]
  reg  valid_144; // @[Icache.scala 18:24]
  reg  valid_145; // @[Icache.scala 18:24]
  reg  valid_146; // @[Icache.scala 18:24]
  reg  valid_147; // @[Icache.scala 18:24]
  reg  valid_148; // @[Icache.scala 18:24]
  reg  valid_149; // @[Icache.scala 18:24]
  reg  valid_150; // @[Icache.scala 18:24]
  reg  valid_151; // @[Icache.scala 18:24]
  reg  valid_152; // @[Icache.scala 18:24]
  reg  valid_153; // @[Icache.scala 18:24]
  reg  valid_154; // @[Icache.scala 18:24]
  reg  valid_155; // @[Icache.scala 18:24]
  reg  valid_156; // @[Icache.scala 18:24]
  reg  valid_157; // @[Icache.scala 18:24]
  reg  valid_158; // @[Icache.scala 18:24]
  reg  valid_159; // @[Icache.scala 18:24]
  reg  valid_160; // @[Icache.scala 18:24]
  reg  valid_161; // @[Icache.scala 18:24]
  reg  valid_162; // @[Icache.scala 18:24]
  reg  valid_163; // @[Icache.scala 18:24]
  reg  valid_164; // @[Icache.scala 18:24]
  reg  valid_165; // @[Icache.scala 18:24]
  reg  valid_166; // @[Icache.scala 18:24]
  reg  valid_167; // @[Icache.scala 18:24]
  reg  valid_168; // @[Icache.scala 18:24]
  reg  valid_169; // @[Icache.scala 18:24]
  reg  valid_170; // @[Icache.scala 18:24]
  reg  valid_171; // @[Icache.scala 18:24]
  reg  valid_172; // @[Icache.scala 18:24]
  reg  valid_173; // @[Icache.scala 18:24]
  reg  valid_174; // @[Icache.scala 18:24]
  reg  valid_175; // @[Icache.scala 18:24]
  reg  valid_176; // @[Icache.scala 18:24]
  reg  valid_177; // @[Icache.scala 18:24]
  reg  valid_178; // @[Icache.scala 18:24]
  reg  valid_179; // @[Icache.scala 18:24]
  reg  valid_180; // @[Icache.scala 18:24]
  reg  valid_181; // @[Icache.scala 18:24]
  reg  valid_182; // @[Icache.scala 18:24]
  reg  valid_183; // @[Icache.scala 18:24]
  reg  valid_184; // @[Icache.scala 18:24]
  reg  valid_185; // @[Icache.scala 18:24]
  reg  valid_186; // @[Icache.scala 18:24]
  reg  valid_187; // @[Icache.scala 18:24]
  reg  valid_188; // @[Icache.scala 18:24]
  reg  valid_189; // @[Icache.scala 18:24]
  reg  valid_190; // @[Icache.scala 18:24]
  reg  valid_191; // @[Icache.scala 18:24]
  reg  valid_192; // @[Icache.scala 18:24]
  reg  valid_193; // @[Icache.scala 18:24]
  reg  valid_194; // @[Icache.scala 18:24]
  reg  valid_195; // @[Icache.scala 18:24]
  reg  valid_196; // @[Icache.scala 18:24]
  reg  valid_197; // @[Icache.scala 18:24]
  reg  valid_198; // @[Icache.scala 18:24]
  reg  valid_199; // @[Icache.scala 18:24]
  reg  valid_200; // @[Icache.scala 18:24]
  reg  valid_201; // @[Icache.scala 18:24]
  reg  valid_202; // @[Icache.scala 18:24]
  reg  valid_203; // @[Icache.scala 18:24]
  reg  valid_204; // @[Icache.scala 18:24]
  reg  valid_205; // @[Icache.scala 18:24]
  reg  valid_206; // @[Icache.scala 18:24]
  reg  valid_207; // @[Icache.scala 18:24]
  reg  valid_208; // @[Icache.scala 18:24]
  reg  valid_209; // @[Icache.scala 18:24]
  reg  valid_210; // @[Icache.scala 18:24]
  reg  valid_211; // @[Icache.scala 18:24]
  reg  valid_212; // @[Icache.scala 18:24]
  reg  valid_213; // @[Icache.scala 18:24]
  reg  valid_214; // @[Icache.scala 18:24]
  reg  valid_215; // @[Icache.scala 18:24]
  reg  valid_216; // @[Icache.scala 18:24]
  reg  valid_217; // @[Icache.scala 18:24]
  reg  valid_218; // @[Icache.scala 18:24]
  reg  valid_219; // @[Icache.scala 18:24]
  reg  valid_220; // @[Icache.scala 18:24]
  reg  valid_221; // @[Icache.scala 18:24]
  reg  valid_222; // @[Icache.scala 18:24]
  reg  valid_223; // @[Icache.scala 18:24]
  reg  valid_224; // @[Icache.scala 18:24]
  reg  valid_225; // @[Icache.scala 18:24]
  reg  valid_226; // @[Icache.scala 18:24]
  reg  valid_227; // @[Icache.scala 18:24]
  reg  valid_228; // @[Icache.scala 18:24]
  reg  valid_229; // @[Icache.scala 18:24]
  reg  valid_230; // @[Icache.scala 18:24]
  reg  valid_231; // @[Icache.scala 18:24]
  reg  valid_232; // @[Icache.scala 18:24]
  reg  valid_233; // @[Icache.scala 18:24]
  reg  valid_234; // @[Icache.scala 18:24]
  reg  valid_235; // @[Icache.scala 18:24]
  reg  valid_236; // @[Icache.scala 18:24]
  reg  valid_237; // @[Icache.scala 18:24]
  reg  valid_238; // @[Icache.scala 18:24]
  reg  valid_239; // @[Icache.scala 18:24]
  reg  valid_240; // @[Icache.scala 18:24]
  reg  valid_241; // @[Icache.scala 18:24]
  reg  valid_242; // @[Icache.scala 18:24]
  reg  valid_243; // @[Icache.scala 18:24]
  reg  valid_244; // @[Icache.scala 18:24]
  reg  valid_245; // @[Icache.scala 18:24]
  reg  valid_246; // @[Icache.scala 18:24]
  reg  valid_247; // @[Icache.scala 18:24]
  reg  valid_248; // @[Icache.scala 18:24]
  reg  valid_249; // @[Icache.scala 18:24]
  reg  valid_250; // @[Icache.scala 18:24]
  reg  valid_251; // @[Icache.scala 18:24]
  reg  valid_252; // @[Icache.scala 18:24]
  reg  valid_253; // @[Icache.scala 18:24]
  reg  valid_254; // @[Icache.scala 18:24]
  reg  valid_255; // @[Icache.scala 18:24]
  reg [2:0] state; // @[Icache.scala 26:22]
  wire [19:0] req_tag = io_imem_inst_addr[31:12]; // @[Icache.scala 28:30]
  wire [7:0] req_index = io_imem_inst_addr[11:4]; // @[Icache.scala 29:30]
  wire [3:0] req_offset = io_imem_inst_addr[3:0]; // @[Icache.scala 30:30]
  wire [19:0] _GEN_1 = 8'h1 == req_index ? tag_1 : tag_0; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_2 = 8'h2 == req_index ? tag_2 : _GEN_1; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_3 = 8'h3 == req_index ? tag_3 : _GEN_2; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_4 = 8'h4 == req_index ? tag_4 : _GEN_3; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_5 = 8'h5 == req_index ? tag_5 : _GEN_4; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_6 = 8'h6 == req_index ? tag_6 : _GEN_5; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_7 = 8'h7 == req_index ? tag_7 : _GEN_6; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_8 = 8'h8 == req_index ? tag_8 : _GEN_7; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_9 = 8'h9 == req_index ? tag_9 : _GEN_8; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_10 = 8'ha == req_index ? tag_10 : _GEN_9; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_11 = 8'hb == req_index ? tag_11 : _GEN_10; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_12 = 8'hc == req_index ? tag_12 : _GEN_11; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_13 = 8'hd == req_index ? tag_13 : _GEN_12; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_14 = 8'he == req_index ? tag_14 : _GEN_13; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_15 = 8'hf == req_index ? tag_15 : _GEN_14; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_16 = 8'h10 == req_index ? tag_16 : _GEN_15; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_17 = 8'h11 == req_index ? tag_17 : _GEN_16; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_18 = 8'h12 == req_index ? tag_18 : _GEN_17; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_19 = 8'h13 == req_index ? tag_19 : _GEN_18; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_20 = 8'h14 == req_index ? tag_20 : _GEN_19; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_21 = 8'h15 == req_index ? tag_21 : _GEN_20; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_22 = 8'h16 == req_index ? tag_22 : _GEN_21; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_23 = 8'h17 == req_index ? tag_23 : _GEN_22; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_24 = 8'h18 == req_index ? tag_24 : _GEN_23; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_25 = 8'h19 == req_index ? tag_25 : _GEN_24; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_26 = 8'h1a == req_index ? tag_26 : _GEN_25; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_27 = 8'h1b == req_index ? tag_27 : _GEN_26; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_28 = 8'h1c == req_index ? tag_28 : _GEN_27; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_29 = 8'h1d == req_index ? tag_29 : _GEN_28; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_30 = 8'h1e == req_index ? tag_30 : _GEN_29; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_31 = 8'h1f == req_index ? tag_31 : _GEN_30; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_32 = 8'h20 == req_index ? tag_32 : _GEN_31; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_33 = 8'h21 == req_index ? tag_33 : _GEN_32; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_34 = 8'h22 == req_index ? tag_34 : _GEN_33; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_35 = 8'h23 == req_index ? tag_35 : _GEN_34; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_36 = 8'h24 == req_index ? tag_36 : _GEN_35; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_37 = 8'h25 == req_index ? tag_37 : _GEN_36; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_38 = 8'h26 == req_index ? tag_38 : _GEN_37; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_39 = 8'h27 == req_index ? tag_39 : _GEN_38; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_40 = 8'h28 == req_index ? tag_40 : _GEN_39; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_41 = 8'h29 == req_index ? tag_41 : _GEN_40; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_42 = 8'h2a == req_index ? tag_42 : _GEN_41; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_43 = 8'h2b == req_index ? tag_43 : _GEN_42; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_44 = 8'h2c == req_index ? tag_44 : _GEN_43; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_45 = 8'h2d == req_index ? tag_45 : _GEN_44; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_46 = 8'h2e == req_index ? tag_46 : _GEN_45; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_47 = 8'h2f == req_index ? tag_47 : _GEN_46; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_48 = 8'h30 == req_index ? tag_48 : _GEN_47; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_49 = 8'h31 == req_index ? tag_49 : _GEN_48; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_50 = 8'h32 == req_index ? tag_50 : _GEN_49; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_51 = 8'h33 == req_index ? tag_51 : _GEN_50; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_52 = 8'h34 == req_index ? tag_52 : _GEN_51; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_53 = 8'h35 == req_index ? tag_53 : _GEN_52; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_54 = 8'h36 == req_index ? tag_54 : _GEN_53; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_55 = 8'h37 == req_index ? tag_55 : _GEN_54; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_56 = 8'h38 == req_index ? tag_56 : _GEN_55; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_57 = 8'h39 == req_index ? tag_57 : _GEN_56; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_58 = 8'h3a == req_index ? tag_58 : _GEN_57; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_59 = 8'h3b == req_index ? tag_59 : _GEN_58; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_60 = 8'h3c == req_index ? tag_60 : _GEN_59; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_61 = 8'h3d == req_index ? tag_61 : _GEN_60; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_62 = 8'h3e == req_index ? tag_62 : _GEN_61; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_63 = 8'h3f == req_index ? tag_63 : _GEN_62; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_64 = 8'h40 == req_index ? tag_64 : _GEN_63; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_65 = 8'h41 == req_index ? tag_65 : _GEN_64; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_66 = 8'h42 == req_index ? tag_66 : _GEN_65; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_67 = 8'h43 == req_index ? tag_67 : _GEN_66; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_68 = 8'h44 == req_index ? tag_68 : _GEN_67; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_69 = 8'h45 == req_index ? tag_69 : _GEN_68; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_70 = 8'h46 == req_index ? tag_70 : _GEN_69; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_71 = 8'h47 == req_index ? tag_71 : _GEN_70; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_72 = 8'h48 == req_index ? tag_72 : _GEN_71; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_73 = 8'h49 == req_index ? tag_73 : _GEN_72; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_74 = 8'h4a == req_index ? tag_74 : _GEN_73; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_75 = 8'h4b == req_index ? tag_75 : _GEN_74; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_76 = 8'h4c == req_index ? tag_76 : _GEN_75; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_77 = 8'h4d == req_index ? tag_77 : _GEN_76; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_78 = 8'h4e == req_index ? tag_78 : _GEN_77; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_79 = 8'h4f == req_index ? tag_79 : _GEN_78; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_80 = 8'h50 == req_index ? tag_80 : _GEN_79; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_81 = 8'h51 == req_index ? tag_81 : _GEN_80; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_82 = 8'h52 == req_index ? tag_82 : _GEN_81; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_83 = 8'h53 == req_index ? tag_83 : _GEN_82; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_84 = 8'h54 == req_index ? tag_84 : _GEN_83; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_85 = 8'h55 == req_index ? tag_85 : _GEN_84; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_86 = 8'h56 == req_index ? tag_86 : _GEN_85; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_87 = 8'h57 == req_index ? tag_87 : _GEN_86; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_88 = 8'h58 == req_index ? tag_88 : _GEN_87; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_89 = 8'h59 == req_index ? tag_89 : _GEN_88; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_90 = 8'h5a == req_index ? tag_90 : _GEN_89; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_91 = 8'h5b == req_index ? tag_91 : _GEN_90; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_92 = 8'h5c == req_index ? tag_92 : _GEN_91; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_93 = 8'h5d == req_index ? tag_93 : _GEN_92; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_94 = 8'h5e == req_index ? tag_94 : _GEN_93; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_95 = 8'h5f == req_index ? tag_95 : _GEN_94; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_96 = 8'h60 == req_index ? tag_96 : _GEN_95; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_97 = 8'h61 == req_index ? tag_97 : _GEN_96; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_98 = 8'h62 == req_index ? tag_98 : _GEN_97; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_99 = 8'h63 == req_index ? tag_99 : _GEN_98; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_100 = 8'h64 == req_index ? tag_100 : _GEN_99; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_101 = 8'h65 == req_index ? tag_101 : _GEN_100; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_102 = 8'h66 == req_index ? tag_102 : _GEN_101; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_103 = 8'h67 == req_index ? tag_103 : _GEN_102; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_104 = 8'h68 == req_index ? tag_104 : _GEN_103; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_105 = 8'h69 == req_index ? tag_105 : _GEN_104; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_106 = 8'h6a == req_index ? tag_106 : _GEN_105; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_107 = 8'h6b == req_index ? tag_107 : _GEN_106; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_108 = 8'h6c == req_index ? tag_108 : _GEN_107; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_109 = 8'h6d == req_index ? tag_109 : _GEN_108; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_110 = 8'h6e == req_index ? tag_110 : _GEN_109; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_111 = 8'h6f == req_index ? tag_111 : _GEN_110; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_112 = 8'h70 == req_index ? tag_112 : _GEN_111; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_113 = 8'h71 == req_index ? tag_113 : _GEN_112; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_114 = 8'h72 == req_index ? tag_114 : _GEN_113; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_115 = 8'h73 == req_index ? tag_115 : _GEN_114; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_116 = 8'h74 == req_index ? tag_116 : _GEN_115; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_117 = 8'h75 == req_index ? tag_117 : _GEN_116; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_118 = 8'h76 == req_index ? tag_118 : _GEN_117; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_119 = 8'h77 == req_index ? tag_119 : _GEN_118; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_120 = 8'h78 == req_index ? tag_120 : _GEN_119; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_121 = 8'h79 == req_index ? tag_121 : _GEN_120; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_122 = 8'h7a == req_index ? tag_122 : _GEN_121; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_123 = 8'h7b == req_index ? tag_123 : _GEN_122; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_124 = 8'h7c == req_index ? tag_124 : _GEN_123; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_125 = 8'h7d == req_index ? tag_125 : _GEN_124; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_126 = 8'h7e == req_index ? tag_126 : _GEN_125; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_127 = 8'h7f == req_index ? tag_127 : _GEN_126; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_128 = 8'h80 == req_index ? tag_128 : _GEN_127; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_129 = 8'h81 == req_index ? tag_129 : _GEN_128; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_130 = 8'h82 == req_index ? tag_130 : _GEN_129; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_131 = 8'h83 == req_index ? tag_131 : _GEN_130; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_132 = 8'h84 == req_index ? tag_132 : _GEN_131; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_133 = 8'h85 == req_index ? tag_133 : _GEN_132; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_134 = 8'h86 == req_index ? tag_134 : _GEN_133; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_135 = 8'h87 == req_index ? tag_135 : _GEN_134; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_136 = 8'h88 == req_index ? tag_136 : _GEN_135; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_137 = 8'h89 == req_index ? tag_137 : _GEN_136; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_138 = 8'h8a == req_index ? tag_138 : _GEN_137; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_139 = 8'h8b == req_index ? tag_139 : _GEN_138; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_140 = 8'h8c == req_index ? tag_140 : _GEN_139; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_141 = 8'h8d == req_index ? tag_141 : _GEN_140; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_142 = 8'h8e == req_index ? tag_142 : _GEN_141; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_143 = 8'h8f == req_index ? tag_143 : _GEN_142; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_144 = 8'h90 == req_index ? tag_144 : _GEN_143; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_145 = 8'h91 == req_index ? tag_145 : _GEN_144; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_146 = 8'h92 == req_index ? tag_146 : _GEN_145; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_147 = 8'h93 == req_index ? tag_147 : _GEN_146; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_148 = 8'h94 == req_index ? tag_148 : _GEN_147; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_149 = 8'h95 == req_index ? tag_149 : _GEN_148; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_150 = 8'h96 == req_index ? tag_150 : _GEN_149; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_151 = 8'h97 == req_index ? tag_151 : _GEN_150; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_152 = 8'h98 == req_index ? tag_152 : _GEN_151; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_153 = 8'h99 == req_index ? tag_153 : _GEN_152; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_154 = 8'h9a == req_index ? tag_154 : _GEN_153; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_155 = 8'h9b == req_index ? tag_155 : _GEN_154; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_156 = 8'h9c == req_index ? tag_156 : _GEN_155; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_157 = 8'h9d == req_index ? tag_157 : _GEN_156; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_158 = 8'h9e == req_index ? tag_158 : _GEN_157; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_159 = 8'h9f == req_index ? tag_159 : _GEN_158; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_160 = 8'ha0 == req_index ? tag_160 : _GEN_159; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_161 = 8'ha1 == req_index ? tag_161 : _GEN_160; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_162 = 8'ha2 == req_index ? tag_162 : _GEN_161; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_163 = 8'ha3 == req_index ? tag_163 : _GEN_162; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_164 = 8'ha4 == req_index ? tag_164 : _GEN_163; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_165 = 8'ha5 == req_index ? tag_165 : _GEN_164; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_166 = 8'ha6 == req_index ? tag_166 : _GEN_165; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_167 = 8'ha7 == req_index ? tag_167 : _GEN_166; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_168 = 8'ha8 == req_index ? tag_168 : _GEN_167; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_169 = 8'ha9 == req_index ? tag_169 : _GEN_168; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_170 = 8'haa == req_index ? tag_170 : _GEN_169; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_171 = 8'hab == req_index ? tag_171 : _GEN_170; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_172 = 8'hac == req_index ? tag_172 : _GEN_171; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_173 = 8'had == req_index ? tag_173 : _GEN_172; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_174 = 8'hae == req_index ? tag_174 : _GEN_173; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_175 = 8'haf == req_index ? tag_175 : _GEN_174; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_176 = 8'hb0 == req_index ? tag_176 : _GEN_175; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_177 = 8'hb1 == req_index ? tag_177 : _GEN_176; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_178 = 8'hb2 == req_index ? tag_178 : _GEN_177; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_179 = 8'hb3 == req_index ? tag_179 : _GEN_178; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_180 = 8'hb4 == req_index ? tag_180 : _GEN_179; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_181 = 8'hb5 == req_index ? tag_181 : _GEN_180; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_182 = 8'hb6 == req_index ? tag_182 : _GEN_181; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_183 = 8'hb7 == req_index ? tag_183 : _GEN_182; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_184 = 8'hb8 == req_index ? tag_184 : _GEN_183; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_185 = 8'hb9 == req_index ? tag_185 : _GEN_184; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_186 = 8'hba == req_index ? tag_186 : _GEN_185; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_187 = 8'hbb == req_index ? tag_187 : _GEN_186; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_188 = 8'hbc == req_index ? tag_188 : _GEN_187; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_189 = 8'hbd == req_index ? tag_189 : _GEN_188; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_190 = 8'hbe == req_index ? tag_190 : _GEN_189; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_191 = 8'hbf == req_index ? tag_191 : _GEN_190; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_192 = 8'hc0 == req_index ? tag_192 : _GEN_191; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_193 = 8'hc1 == req_index ? tag_193 : _GEN_192; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_194 = 8'hc2 == req_index ? tag_194 : _GEN_193; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_195 = 8'hc3 == req_index ? tag_195 : _GEN_194; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_196 = 8'hc4 == req_index ? tag_196 : _GEN_195; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_197 = 8'hc5 == req_index ? tag_197 : _GEN_196; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_198 = 8'hc6 == req_index ? tag_198 : _GEN_197; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_199 = 8'hc7 == req_index ? tag_199 : _GEN_198; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_200 = 8'hc8 == req_index ? tag_200 : _GEN_199; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_201 = 8'hc9 == req_index ? tag_201 : _GEN_200; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_202 = 8'hca == req_index ? tag_202 : _GEN_201; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_203 = 8'hcb == req_index ? tag_203 : _GEN_202; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_204 = 8'hcc == req_index ? tag_204 : _GEN_203; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_205 = 8'hcd == req_index ? tag_205 : _GEN_204; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_206 = 8'hce == req_index ? tag_206 : _GEN_205; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_207 = 8'hcf == req_index ? tag_207 : _GEN_206; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_208 = 8'hd0 == req_index ? tag_208 : _GEN_207; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_209 = 8'hd1 == req_index ? tag_209 : _GEN_208; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_210 = 8'hd2 == req_index ? tag_210 : _GEN_209; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_211 = 8'hd3 == req_index ? tag_211 : _GEN_210; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_212 = 8'hd4 == req_index ? tag_212 : _GEN_211; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_213 = 8'hd5 == req_index ? tag_213 : _GEN_212; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_214 = 8'hd6 == req_index ? tag_214 : _GEN_213; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_215 = 8'hd7 == req_index ? tag_215 : _GEN_214; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_216 = 8'hd8 == req_index ? tag_216 : _GEN_215; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_217 = 8'hd9 == req_index ? tag_217 : _GEN_216; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_218 = 8'hda == req_index ? tag_218 : _GEN_217; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_219 = 8'hdb == req_index ? tag_219 : _GEN_218; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_220 = 8'hdc == req_index ? tag_220 : _GEN_219; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_221 = 8'hdd == req_index ? tag_221 : _GEN_220; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_222 = 8'hde == req_index ? tag_222 : _GEN_221; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_223 = 8'hdf == req_index ? tag_223 : _GEN_222; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_224 = 8'he0 == req_index ? tag_224 : _GEN_223; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_225 = 8'he1 == req_index ? tag_225 : _GEN_224; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_226 = 8'he2 == req_index ? tag_226 : _GEN_225; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_227 = 8'he3 == req_index ? tag_227 : _GEN_226; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_228 = 8'he4 == req_index ? tag_228 : _GEN_227; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_229 = 8'he5 == req_index ? tag_229 : _GEN_228; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_230 = 8'he6 == req_index ? tag_230 : _GEN_229; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_231 = 8'he7 == req_index ? tag_231 : _GEN_230; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_232 = 8'he8 == req_index ? tag_232 : _GEN_231; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_233 = 8'he9 == req_index ? tag_233 : _GEN_232; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_234 = 8'hea == req_index ? tag_234 : _GEN_233; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_235 = 8'heb == req_index ? tag_235 : _GEN_234; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_236 = 8'hec == req_index ? tag_236 : _GEN_235; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_237 = 8'hed == req_index ? tag_237 : _GEN_236; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_238 = 8'hee == req_index ? tag_238 : _GEN_237; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_239 = 8'hef == req_index ? tag_239 : _GEN_238; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_240 = 8'hf0 == req_index ? tag_240 : _GEN_239; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_241 = 8'hf1 == req_index ? tag_241 : _GEN_240; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_242 = 8'hf2 == req_index ? tag_242 : _GEN_241; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_243 = 8'hf3 == req_index ? tag_243 : _GEN_242; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_244 = 8'hf4 == req_index ? tag_244 : _GEN_243; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_245 = 8'hf5 == req_index ? tag_245 : _GEN_244; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_246 = 8'hf6 == req_index ? tag_246 : _GEN_245; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_247 = 8'hf7 == req_index ? tag_247 : _GEN_246; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_248 = 8'hf8 == req_index ? tag_248 : _GEN_247; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_249 = 8'hf9 == req_index ? tag_249 : _GEN_248; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_250 = 8'hfa == req_index ? tag_250 : _GEN_249; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_251 = 8'hfb == req_index ? tag_251 : _GEN_250; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_252 = 8'hfc == req_index ? tag_252 : _GEN_251; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_253 = 8'hfd == req_index ? tag_253 : _GEN_252; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_254 = 8'hfe == req_index ? tag_254 : _GEN_253; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire [19:0] _GEN_255 = 8'hff == req_index ? tag_255 : _GEN_254; // @[Icache.scala 33:32 Icache.scala 33:32]
  wire  _GEN_257 = 8'h1 == req_index ? valid_1 : valid_0; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_258 = 8'h2 == req_index ? valid_2 : _GEN_257; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_259 = 8'h3 == req_index ? valid_3 : _GEN_258; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_260 = 8'h4 == req_index ? valid_4 : _GEN_259; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_261 = 8'h5 == req_index ? valid_5 : _GEN_260; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_262 = 8'h6 == req_index ? valid_6 : _GEN_261; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_263 = 8'h7 == req_index ? valid_7 : _GEN_262; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_264 = 8'h8 == req_index ? valid_8 : _GEN_263; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_265 = 8'h9 == req_index ? valid_9 : _GEN_264; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_266 = 8'ha == req_index ? valid_10 : _GEN_265; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_267 = 8'hb == req_index ? valid_11 : _GEN_266; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_268 = 8'hc == req_index ? valid_12 : _GEN_267; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_269 = 8'hd == req_index ? valid_13 : _GEN_268; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_270 = 8'he == req_index ? valid_14 : _GEN_269; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_271 = 8'hf == req_index ? valid_15 : _GEN_270; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_272 = 8'h10 == req_index ? valid_16 : _GEN_271; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_273 = 8'h11 == req_index ? valid_17 : _GEN_272; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_274 = 8'h12 == req_index ? valid_18 : _GEN_273; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_275 = 8'h13 == req_index ? valid_19 : _GEN_274; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_276 = 8'h14 == req_index ? valid_20 : _GEN_275; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_277 = 8'h15 == req_index ? valid_21 : _GEN_276; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_278 = 8'h16 == req_index ? valid_22 : _GEN_277; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_279 = 8'h17 == req_index ? valid_23 : _GEN_278; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_280 = 8'h18 == req_index ? valid_24 : _GEN_279; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_281 = 8'h19 == req_index ? valid_25 : _GEN_280; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_282 = 8'h1a == req_index ? valid_26 : _GEN_281; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_283 = 8'h1b == req_index ? valid_27 : _GEN_282; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_284 = 8'h1c == req_index ? valid_28 : _GEN_283; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_285 = 8'h1d == req_index ? valid_29 : _GEN_284; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_286 = 8'h1e == req_index ? valid_30 : _GEN_285; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_287 = 8'h1f == req_index ? valid_31 : _GEN_286; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_288 = 8'h20 == req_index ? valid_32 : _GEN_287; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_289 = 8'h21 == req_index ? valid_33 : _GEN_288; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_290 = 8'h22 == req_index ? valid_34 : _GEN_289; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_291 = 8'h23 == req_index ? valid_35 : _GEN_290; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_292 = 8'h24 == req_index ? valid_36 : _GEN_291; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_293 = 8'h25 == req_index ? valid_37 : _GEN_292; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_294 = 8'h26 == req_index ? valid_38 : _GEN_293; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_295 = 8'h27 == req_index ? valid_39 : _GEN_294; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_296 = 8'h28 == req_index ? valid_40 : _GEN_295; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_297 = 8'h29 == req_index ? valid_41 : _GEN_296; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_298 = 8'h2a == req_index ? valid_42 : _GEN_297; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_299 = 8'h2b == req_index ? valid_43 : _GEN_298; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_300 = 8'h2c == req_index ? valid_44 : _GEN_299; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_301 = 8'h2d == req_index ? valid_45 : _GEN_300; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_302 = 8'h2e == req_index ? valid_46 : _GEN_301; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_303 = 8'h2f == req_index ? valid_47 : _GEN_302; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_304 = 8'h30 == req_index ? valid_48 : _GEN_303; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_305 = 8'h31 == req_index ? valid_49 : _GEN_304; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_306 = 8'h32 == req_index ? valid_50 : _GEN_305; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_307 = 8'h33 == req_index ? valid_51 : _GEN_306; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_308 = 8'h34 == req_index ? valid_52 : _GEN_307; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_309 = 8'h35 == req_index ? valid_53 : _GEN_308; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_310 = 8'h36 == req_index ? valid_54 : _GEN_309; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_311 = 8'h37 == req_index ? valid_55 : _GEN_310; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_312 = 8'h38 == req_index ? valid_56 : _GEN_311; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_313 = 8'h39 == req_index ? valid_57 : _GEN_312; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_314 = 8'h3a == req_index ? valid_58 : _GEN_313; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_315 = 8'h3b == req_index ? valid_59 : _GEN_314; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_316 = 8'h3c == req_index ? valid_60 : _GEN_315; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_317 = 8'h3d == req_index ? valid_61 : _GEN_316; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_318 = 8'h3e == req_index ? valid_62 : _GEN_317; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_319 = 8'h3f == req_index ? valid_63 : _GEN_318; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_320 = 8'h40 == req_index ? valid_64 : _GEN_319; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_321 = 8'h41 == req_index ? valid_65 : _GEN_320; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_322 = 8'h42 == req_index ? valid_66 : _GEN_321; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_323 = 8'h43 == req_index ? valid_67 : _GEN_322; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_324 = 8'h44 == req_index ? valid_68 : _GEN_323; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_325 = 8'h45 == req_index ? valid_69 : _GEN_324; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_326 = 8'h46 == req_index ? valid_70 : _GEN_325; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_327 = 8'h47 == req_index ? valid_71 : _GEN_326; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_328 = 8'h48 == req_index ? valid_72 : _GEN_327; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_329 = 8'h49 == req_index ? valid_73 : _GEN_328; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_330 = 8'h4a == req_index ? valid_74 : _GEN_329; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_331 = 8'h4b == req_index ? valid_75 : _GEN_330; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_332 = 8'h4c == req_index ? valid_76 : _GEN_331; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_333 = 8'h4d == req_index ? valid_77 : _GEN_332; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_334 = 8'h4e == req_index ? valid_78 : _GEN_333; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_335 = 8'h4f == req_index ? valid_79 : _GEN_334; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_336 = 8'h50 == req_index ? valid_80 : _GEN_335; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_337 = 8'h51 == req_index ? valid_81 : _GEN_336; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_338 = 8'h52 == req_index ? valid_82 : _GEN_337; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_339 = 8'h53 == req_index ? valid_83 : _GEN_338; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_340 = 8'h54 == req_index ? valid_84 : _GEN_339; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_341 = 8'h55 == req_index ? valid_85 : _GEN_340; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_342 = 8'h56 == req_index ? valid_86 : _GEN_341; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_343 = 8'h57 == req_index ? valid_87 : _GEN_342; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_344 = 8'h58 == req_index ? valid_88 : _GEN_343; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_345 = 8'h59 == req_index ? valid_89 : _GEN_344; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_346 = 8'h5a == req_index ? valid_90 : _GEN_345; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_347 = 8'h5b == req_index ? valid_91 : _GEN_346; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_348 = 8'h5c == req_index ? valid_92 : _GEN_347; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_349 = 8'h5d == req_index ? valid_93 : _GEN_348; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_350 = 8'h5e == req_index ? valid_94 : _GEN_349; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_351 = 8'h5f == req_index ? valid_95 : _GEN_350; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_352 = 8'h60 == req_index ? valid_96 : _GEN_351; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_353 = 8'h61 == req_index ? valid_97 : _GEN_352; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_354 = 8'h62 == req_index ? valid_98 : _GEN_353; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_355 = 8'h63 == req_index ? valid_99 : _GEN_354; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_356 = 8'h64 == req_index ? valid_100 : _GEN_355; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_357 = 8'h65 == req_index ? valid_101 : _GEN_356; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_358 = 8'h66 == req_index ? valid_102 : _GEN_357; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_359 = 8'h67 == req_index ? valid_103 : _GEN_358; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_360 = 8'h68 == req_index ? valid_104 : _GEN_359; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_361 = 8'h69 == req_index ? valid_105 : _GEN_360; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_362 = 8'h6a == req_index ? valid_106 : _GEN_361; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_363 = 8'h6b == req_index ? valid_107 : _GEN_362; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_364 = 8'h6c == req_index ? valid_108 : _GEN_363; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_365 = 8'h6d == req_index ? valid_109 : _GEN_364; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_366 = 8'h6e == req_index ? valid_110 : _GEN_365; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_367 = 8'h6f == req_index ? valid_111 : _GEN_366; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_368 = 8'h70 == req_index ? valid_112 : _GEN_367; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_369 = 8'h71 == req_index ? valid_113 : _GEN_368; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_370 = 8'h72 == req_index ? valid_114 : _GEN_369; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_371 = 8'h73 == req_index ? valid_115 : _GEN_370; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_372 = 8'h74 == req_index ? valid_116 : _GEN_371; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_373 = 8'h75 == req_index ? valid_117 : _GEN_372; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_374 = 8'h76 == req_index ? valid_118 : _GEN_373; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_375 = 8'h77 == req_index ? valid_119 : _GEN_374; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_376 = 8'h78 == req_index ? valid_120 : _GEN_375; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_377 = 8'h79 == req_index ? valid_121 : _GEN_376; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_378 = 8'h7a == req_index ? valid_122 : _GEN_377; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_379 = 8'h7b == req_index ? valid_123 : _GEN_378; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_380 = 8'h7c == req_index ? valid_124 : _GEN_379; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_381 = 8'h7d == req_index ? valid_125 : _GEN_380; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_382 = 8'h7e == req_index ? valid_126 : _GEN_381; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_383 = 8'h7f == req_index ? valid_127 : _GEN_382; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_384 = 8'h80 == req_index ? valid_128 : _GEN_383; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_385 = 8'h81 == req_index ? valid_129 : _GEN_384; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_386 = 8'h82 == req_index ? valid_130 : _GEN_385; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_387 = 8'h83 == req_index ? valid_131 : _GEN_386; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_388 = 8'h84 == req_index ? valid_132 : _GEN_387; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_389 = 8'h85 == req_index ? valid_133 : _GEN_388; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_390 = 8'h86 == req_index ? valid_134 : _GEN_389; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_391 = 8'h87 == req_index ? valid_135 : _GEN_390; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_392 = 8'h88 == req_index ? valid_136 : _GEN_391; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_393 = 8'h89 == req_index ? valid_137 : _GEN_392; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_394 = 8'h8a == req_index ? valid_138 : _GEN_393; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_395 = 8'h8b == req_index ? valid_139 : _GEN_394; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_396 = 8'h8c == req_index ? valid_140 : _GEN_395; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_397 = 8'h8d == req_index ? valid_141 : _GEN_396; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_398 = 8'h8e == req_index ? valid_142 : _GEN_397; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_399 = 8'h8f == req_index ? valid_143 : _GEN_398; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_400 = 8'h90 == req_index ? valid_144 : _GEN_399; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_401 = 8'h91 == req_index ? valid_145 : _GEN_400; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_402 = 8'h92 == req_index ? valid_146 : _GEN_401; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_403 = 8'h93 == req_index ? valid_147 : _GEN_402; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_404 = 8'h94 == req_index ? valid_148 : _GEN_403; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_405 = 8'h95 == req_index ? valid_149 : _GEN_404; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_406 = 8'h96 == req_index ? valid_150 : _GEN_405; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_407 = 8'h97 == req_index ? valid_151 : _GEN_406; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_408 = 8'h98 == req_index ? valid_152 : _GEN_407; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_409 = 8'h99 == req_index ? valid_153 : _GEN_408; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_410 = 8'h9a == req_index ? valid_154 : _GEN_409; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_411 = 8'h9b == req_index ? valid_155 : _GEN_410; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_412 = 8'h9c == req_index ? valid_156 : _GEN_411; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_413 = 8'h9d == req_index ? valid_157 : _GEN_412; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_414 = 8'h9e == req_index ? valid_158 : _GEN_413; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_415 = 8'h9f == req_index ? valid_159 : _GEN_414; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_416 = 8'ha0 == req_index ? valid_160 : _GEN_415; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_417 = 8'ha1 == req_index ? valid_161 : _GEN_416; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_418 = 8'ha2 == req_index ? valid_162 : _GEN_417; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_419 = 8'ha3 == req_index ? valid_163 : _GEN_418; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_420 = 8'ha4 == req_index ? valid_164 : _GEN_419; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_421 = 8'ha5 == req_index ? valid_165 : _GEN_420; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_422 = 8'ha6 == req_index ? valid_166 : _GEN_421; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_423 = 8'ha7 == req_index ? valid_167 : _GEN_422; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_424 = 8'ha8 == req_index ? valid_168 : _GEN_423; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_425 = 8'ha9 == req_index ? valid_169 : _GEN_424; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_426 = 8'haa == req_index ? valid_170 : _GEN_425; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_427 = 8'hab == req_index ? valid_171 : _GEN_426; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_428 = 8'hac == req_index ? valid_172 : _GEN_427; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_429 = 8'had == req_index ? valid_173 : _GEN_428; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_430 = 8'hae == req_index ? valid_174 : _GEN_429; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_431 = 8'haf == req_index ? valid_175 : _GEN_430; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_432 = 8'hb0 == req_index ? valid_176 : _GEN_431; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_433 = 8'hb1 == req_index ? valid_177 : _GEN_432; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_434 = 8'hb2 == req_index ? valid_178 : _GEN_433; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_435 = 8'hb3 == req_index ? valid_179 : _GEN_434; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_436 = 8'hb4 == req_index ? valid_180 : _GEN_435; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_437 = 8'hb5 == req_index ? valid_181 : _GEN_436; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_438 = 8'hb6 == req_index ? valid_182 : _GEN_437; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_439 = 8'hb7 == req_index ? valid_183 : _GEN_438; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_440 = 8'hb8 == req_index ? valid_184 : _GEN_439; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_441 = 8'hb9 == req_index ? valid_185 : _GEN_440; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_442 = 8'hba == req_index ? valid_186 : _GEN_441; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_443 = 8'hbb == req_index ? valid_187 : _GEN_442; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_444 = 8'hbc == req_index ? valid_188 : _GEN_443; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_445 = 8'hbd == req_index ? valid_189 : _GEN_444; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_446 = 8'hbe == req_index ? valid_190 : _GEN_445; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_447 = 8'hbf == req_index ? valid_191 : _GEN_446; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_448 = 8'hc0 == req_index ? valid_192 : _GEN_447; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_449 = 8'hc1 == req_index ? valid_193 : _GEN_448; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_450 = 8'hc2 == req_index ? valid_194 : _GEN_449; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_451 = 8'hc3 == req_index ? valid_195 : _GEN_450; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_452 = 8'hc4 == req_index ? valid_196 : _GEN_451; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_453 = 8'hc5 == req_index ? valid_197 : _GEN_452; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_454 = 8'hc6 == req_index ? valid_198 : _GEN_453; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_455 = 8'hc7 == req_index ? valid_199 : _GEN_454; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_456 = 8'hc8 == req_index ? valid_200 : _GEN_455; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_457 = 8'hc9 == req_index ? valid_201 : _GEN_456; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_458 = 8'hca == req_index ? valid_202 : _GEN_457; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_459 = 8'hcb == req_index ? valid_203 : _GEN_458; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_460 = 8'hcc == req_index ? valid_204 : _GEN_459; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_461 = 8'hcd == req_index ? valid_205 : _GEN_460; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_462 = 8'hce == req_index ? valid_206 : _GEN_461; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_463 = 8'hcf == req_index ? valid_207 : _GEN_462; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_464 = 8'hd0 == req_index ? valid_208 : _GEN_463; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_465 = 8'hd1 == req_index ? valid_209 : _GEN_464; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_466 = 8'hd2 == req_index ? valid_210 : _GEN_465; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_467 = 8'hd3 == req_index ? valid_211 : _GEN_466; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_468 = 8'hd4 == req_index ? valid_212 : _GEN_467; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_469 = 8'hd5 == req_index ? valid_213 : _GEN_468; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_470 = 8'hd6 == req_index ? valid_214 : _GEN_469; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_471 = 8'hd7 == req_index ? valid_215 : _GEN_470; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_472 = 8'hd8 == req_index ? valid_216 : _GEN_471; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_473 = 8'hd9 == req_index ? valid_217 : _GEN_472; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_474 = 8'hda == req_index ? valid_218 : _GEN_473; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_475 = 8'hdb == req_index ? valid_219 : _GEN_474; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_476 = 8'hdc == req_index ? valid_220 : _GEN_475; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_477 = 8'hdd == req_index ? valid_221 : _GEN_476; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_478 = 8'hde == req_index ? valid_222 : _GEN_477; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_479 = 8'hdf == req_index ? valid_223 : _GEN_478; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_480 = 8'he0 == req_index ? valid_224 : _GEN_479; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_481 = 8'he1 == req_index ? valid_225 : _GEN_480; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_482 = 8'he2 == req_index ? valid_226 : _GEN_481; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_483 = 8'he3 == req_index ? valid_227 : _GEN_482; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_484 = 8'he4 == req_index ? valid_228 : _GEN_483; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_485 = 8'he5 == req_index ? valid_229 : _GEN_484; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_486 = 8'he6 == req_index ? valid_230 : _GEN_485; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_487 = 8'he7 == req_index ? valid_231 : _GEN_486; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_488 = 8'he8 == req_index ? valid_232 : _GEN_487; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_489 = 8'he9 == req_index ? valid_233 : _GEN_488; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_490 = 8'hea == req_index ? valid_234 : _GEN_489; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_491 = 8'heb == req_index ? valid_235 : _GEN_490; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_492 = 8'hec == req_index ? valid_236 : _GEN_491; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_493 = 8'hed == req_index ? valid_237 : _GEN_492; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_494 = 8'hee == req_index ? valid_238 : _GEN_493; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_495 = 8'hef == req_index ? valid_239 : _GEN_494; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_496 = 8'hf0 == req_index ? valid_240 : _GEN_495; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_497 = 8'hf1 == req_index ? valid_241 : _GEN_496; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_498 = 8'hf2 == req_index ? valid_242 : _GEN_497; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_499 = 8'hf3 == req_index ? valid_243 : _GEN_498; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_500 = 8'hf4 == req_index ? valid_244 : _GEN_499; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_501 = 8'hf5 == req_index ? valid_245 : _GEN_500; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_502 = 8'hf6 == req_index ? valid_246 : _GEN_501; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_503 = 8'hf7 == req_index ? valid_247 : _GEN_502; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_504 = 8'hf8 == req_index ? valid_248 : _GEN_503; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_505 = 8'hf9 == req_index ? valid_249 : _GEN_504; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_506 = 8'hfa == req_index ? valid_250 : _GEN_505; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_507 = 8'hfb == req_index ? valid_251 : _GEN_506; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_508 = 8'hfc == req_index ? valid_252 : _GEN_507; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_509 = 8'hfd == req_index ? valid_253 : _GEN_508; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_510 = 8'hfe == req_index ? valid_254 : _GEN_509; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  _GEN_511 = 8'hff == req_index ? valid_255 : _GEN_510; // @[Icache.scala 33:45 Icache.scala 33:45]
  wire  cache_hit = _GEN_255 == req_tag & _GEN_511; // @[Icache.scala 33:45]
  reg  inst_ready; // @[Icache.scala 42:28]
  wire [127:0] cache_data_out = req_Q; // @[Icache.scala 35:28 Icache.scala 132:18]
  wire [31:0] _inst_read_T_6 = 2'h1 == req_offset[3:2] ? cache_data_out[63:32] : cache_data_out[31:0]; // @[Mux.scala 80:57]
  wire [31:0] _inst_read_T_8 = 2'h2 == req_offset[3:2] ? cache_data_out[95:64] : _inst_read_T_6; // @[Mux.scala 80:57]
  reg  cache_fill; // @[Icache.scala 51:28]
  reg  cache_wen; // @[Icache.scala 52:28]
  reg [127:0] cache_wdata; // @[Icache.scala 53:28]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_2 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _GEN_514 = 8'h0 == req_index | valid_0; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_515 = 8'h1 == req_index | valid_1; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_516 = 8'h2 == req_index | valid_2; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_517 = 8'h3 == req_index | valid_3; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_518 = 8'h4 == req_index | valid_4; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_519 = 8'h5 == req_index | valid_5; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_520 = 8'h6 == req_index | valid_6; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_521 = 8'h7 == req_index | valid_7; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_522 = 8'h8 == req_index | valid_8; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_523 = 8'h9 == req_index | valid_9; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_524 = 8'ha == req_index | valid_10; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_525 = 8'hb == req_index | valid_11; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_526 = 8'hc == req_index | valid_12; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_527 = 8'hd == req_index | valid_13; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_528 = 8'he == req_index | valid_14; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_529 = 8'hf == req_index | valid_15; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_530 = 8'h10 == req_index | valid_16; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_531 = 8'h11 == req_index | valid_17; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_532 = 8'h12 == req_index | valid_18; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_533 = 8'h13 == req_index | valid_19; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_534 = 8'h14 == req_index | valid_20; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_535 = 8'h15 == req_index | valid_21; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_536 = 8'h16 == req_index | valid_22; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_537 = 8'h17 == req_index | valid_23; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_538 = 8'h18 == req_index | valid_24; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_539 = 8'h19 == req_index | valid_25; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_540 = 8'h1a == req_index | valid_26; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_541 = 8'h1b == req_index | valid_27; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_542 = 8'h1c == req_index | valid_28; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_543 = 8'h1d == req_index | valid_29; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_544 = 8'h1e == req_index | valid_30; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_545 = 8'h1f == req_index | valid_31; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_546 = 8'h20 == req_index | valid_32; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_547 = 8'h21 == req_index | valid_33; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_548 = 8'h22 == req_index | valid_34; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_549 = 8'h23 == req_index | valid_35; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_550 = 8'h24 == req_index | valid_36; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_551 = 8'h25 == req_index | valid_37; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_552 = 8'h26 == req_index | valid_38; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_553 = 8'h27 == req_index | valid_39; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_554 = 8'h28 == req_index | valid_40; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_555 = 8'h29 == req_index | valid_41; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_556 = 8'h2a == req_index | valid_42; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_557 = 8'h2b == req_index | valid_43; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_558 = 8'h2c == req_index | valid_44; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_559 = 8'h2d == req_index | valid_45; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_560 = 8'h2e == req_index | valid_46; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_561 = 8'h2f == req_index | valid_47; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_562 = 8'h30 == req_index | valid_48; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_563 = 8'h31 == req_index | valid_49; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_564 = 8'h32 == req_index | valid_50; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_565 = 8'h33 == req_index | valid_51; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_566 = 8'h34 == req_index | valid_52; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_567 = 8'h35 == req_index | valid_53; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_568 = 8'h36 == req_index | valid_54; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_569 = 8'h37 == req_index | valid_55; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_570 = 8'h38 == req_index | valid_56; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_571 = 8'h39 == req_index | valid_57; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_572 = 8'h3a == req_index | valid_58; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_573 = 8'h3b == req_index | valid_59; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_574 = 8'h3c == req_index | valid_60; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_575 = 8'h3d == req_index | valid_61; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_576 = 8'h3e == req_index | valid_62; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_577 = 8'h3f == req_index | valid_63; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_578 = 8'h40 == req_index | valid_64; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_579 = 8'h41 == req_index | valid_65; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_580 = 8'h42 == req_index | valid_66; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_581 = 8'h43 == req_index | valid_67; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_582 = 8'h44 == req_index | valid_68; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_583 = 8'h45 == req_index | valid_69; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_584 = 8'h46 == req_index | valid_70; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_585 = 8'h47 == req_index | valid_71; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_586 = 8'h48 == req_index | valid_72; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_587 = 8'h49 == req_index | valid_73; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_588 = 8'h4a == req_index | valid_74; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_589 = 8'h4b == req_index | valid_75; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_590 = 8'h4c == req_index | valid_76; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_591 = 8'h4d == req_index | valid_77; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_592 = 8'h4e == req_index | valid_78; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_593 = 8'h4f == req_index | valid_79; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_594 = 8'h50 == req_index | valid_80; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_595 = 8'h51 == req_index | valid_81; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_596 = 8'h52 == req_index | valid_82; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_597 = 8'h53 == req_index | valid_83; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_598 = 8'h54 == req_index | valid_84; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_599 = 8'h55 == req_index | valid_85; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_600 = 8'h56 == req_index | valid_86; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_601 = 8'h57 == req_index | valid_87; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_602 = 8'h58 == req_index | valid_88; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_603 = 8'h59 == req_index | valid_89; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_604 = 8'h5a == req_index | valid_90; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_605 = 8'h5b == req_index | valid_91; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_606 = 8'h5c == req_index | valid_92; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_607 = 8'h5d == req_index | valid_93; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_608 = 8'h5e == req_index | valid_94; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_609 = 8'h5f == req_index | valid_95; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_610 = 8'h60 == req_index | valid_96; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_611 = 8'h61 == req_index | valid_97; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_612 = 8'h62 == req_index | valid_98; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_613 = 8'h63 == req_index | valid_99; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_614 = 8'h64 == req_index | valid_100; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_615 = 8'h65 == req_index | valid_101; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_616 = 8'h66 == req_index | valid_102; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_617 = 8'h67 == req_index | valid_103; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_618 = 8'h68 == req_index | valid_104; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_619 = 8'h69 == req_index | valid_105; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_620 = 8'h6a == req_index | valid_106; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_621 = 8'h6b == req_index | valid_107; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_622 = 8'h6c == req_index | valid_108; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_623 = 8'h6d == req_index | valid_109; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_624 = 8'h6e == req_index | valid_110; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_625 = 8'h6f == req_index | valid_111; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_626 = 8'h70 == req_index | valid_112; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_627 = 8'h71 == req_index | valid_113; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_628 = 8'h72 == req_index | valid_114; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_629 = 8'h73 == req_index | valid_115; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_630 = 8'h74 == req_index | valid_116; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_631 = 8'h75 == req_index | valid_117; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_632 = 8'h76 == req_index | valid_118; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_633 = 8'h77 == req_index | valid_119; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_634 = 8'h78 == req_index | valid_120; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_635 = 8'h79 == req_index | valid_121; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_636 = 8'h7a == req_index | valid_122; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_637 = 8'h7b == req_index | valid_123; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_638 = 8'h7c == req_index | valid_124; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_639 = 8'h7d == req_index | valid_125; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_640 = 8'h7e == req_index | valid_126; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_641 = 8'h7f == req_index | valid_127; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_642 = 8'h80 == req_index | valid_128; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_643 = 8'h81 == req_index | valid_129; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_644 = 8'h82 == req_index | valid_130; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_645 = 8'h83 == req_index | valid_131; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_646 = 8'h84 == req_index | valid_132; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_647 = 8'h85 == req_index | valid_133; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_648 = 8'h86 == req_index | valid_134; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_649 = 8'h87 == req_index | valid_135; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_650 = 8'h88 == req_index | valid_136; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_651 = 8'h89 == req_index | valid_137; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_652 = 8'h8a == req_index | valid_138; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_653 = 8'h8b == req_index | valid_139; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_654 = 8'h8c == req_index | valid_140; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_655 = 8'h8d == req_index | valid_141; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_656 = 8'h8e == req_index | valid_142; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_657 = 8'h8f == req_index | valid_143; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_658 = 8'h90 == req_index | valid_144; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_659 = 8'h91 == req_index | valid_145; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_660 = 8'h92 == req_index | valid_146; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_661 = 8'h93 == req_index | valid_147; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_662 = 8'h94 == req_index | valid_148; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_663 = 8'h95 == req_index | valid_149; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_664 = 8'h96 == req_index | valid_150; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_665 = 8'h97 == req_index | valid_151; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_666 = 8'h98 == req_index | valid_152; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_667 = 8'h99 == req_index | valid_153; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_668 = 8'h9a == req_index | valid_154; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_669 = 8'h9b == req_index | valid_155; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_670 = 8'h9c == req_index | valid_156; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_671 = 8'h9d == req_index | valid_157; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_672 = 8'h9e == req_index | valid_158; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_673 = 8'h9f == req_index | valid_159; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_674 = 8'ha0 == req_index | valid_160; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_675 = 8'ha1 == req_index | valid_161; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_676 = 8'ha2 == req_index | valid_162; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_677 = 8'ha3 == req_index | valid_163; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_678 = 8'ha4 == req_index | valid_164; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_679 = 8'ha5 == req_index | valid_165; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_680 = 8'ha6 == req_index | valid_166; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_681 = 8'ha7 == req_index | valid_167; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_682 = 8'ha8 == req_index | valid_168; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_683 = 8'ha9 == req_index | valid_169; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_684 = 8'haa == req_index | valid_170; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_685 = 8'hab == req_index | valid_171; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_686 = 8'hac == req_index | valid_172; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_687 = 8'had == req_index | valid_173; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_688 = 8'hae == req_index | valid_174; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_689 = 8'haf == req_index | valid_175; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_690 = 8'hb0 == req_index | valid_176; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_691 = 8'hb1 == req_index | valid_177; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_692 = 8'hb2 == req_index | valid_178; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_693 = 8'hb3 == req_index | valid_179; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_694 = 8'hb4 == req_index | valid_180; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_695 = 8'hb5 == req_index | valid_181; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_696 = 8'hb6 == req_index | valid_182; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_697 = 8'hb7 == req_index | valid_183; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_698 = 8'hb8 == req_index | valid_184; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_699 = 8'hb9 == req_index | valid_185; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_700 = 8'hba == req_index | valid_186; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_701 = 8'hbb == req_index | valid_187; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_702 = 8'hbc == req_index | valid_188; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_703 = 8'hbd == req_index | valid_189; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_704 = 8'hbe == req_index | valid_190; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_705 = 8'hbf == req_index | valid_191; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_706 = 8'hc0 == req_index | valid_192; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_707 = 8'hc1 == req_index | valid_193; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_708 = 8'hc2 == req_index | valid_194; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_709 = 8'hc3 == req_index | valid_195; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_710 = 8'hc4 == req_index | valid_196; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_711 = 8'hc5 == req_index | valid_197; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_712 = 8'hc6 == req_index | valid_198; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_713 = 8'hc7 == req_index | valid_199; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_714 = 8'hc8 == req_index | valid_200; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_715 = 8'hc9 == req_index | valid_201; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_716 = 8'hca == req_index | valid_202; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_717 = 8'hcb == req_index | valid_203; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_718 = 8'hcc == req_index | valid_204; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_719 = 8'hcd == req_index | valid_205; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_720 = 8'hce == req_index | valid_206; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_721 = 8'hcf == req_index | valid_207; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_722 = 8'hd0 == req_index | valid_208; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_723 = 8'hd1 == req_index | valid_209; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_724 = 8'hd2 == req_index | valid_210; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_725 = 8'hd3 == req_index | valid_211; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_726 = 8'hd4 == req_index | valid_212; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_727 = 8'hd5 == req_index | valid_213; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_728 = 8'hd6 == req_index | valid_214; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_729 = 8'hd7 == req_index | valid_215; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_730 = 8'hd8 == req_index | valid_216; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_731 = 8'hd9 == req_index | valid_217; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_732 = 8'hda == req_index | valid_218; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_733 = 8'hdb == req_index | valid_219; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_734 = 8'hdc == req_index | valid_220; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_735 = 8'hdd == req_index | valid_221; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_736 = 8'hde == req_index | valid_222; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_737 = 8'hdf == req_index | valid_223; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_738 = 8'he0 == req_index | valid_224; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_739 = 8'he1 == req_index | valid_225; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_740 = 8'he2 == req_index | valid_226; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_741 = 8'he3 == req_index | valid_227; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_742 = 8'he4 == req_index | valid_228; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_743 = 8'he5 == req_index | valid_229; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_744 = 8'he6 == req_index | valid_230; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_745 = 8'he7 == req_index | valid_231; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_746 = 8'he8 == req_index | valid_232; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_747 = 8'he9 == req_index | valid_233; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_748 = 8'hea == req_index | valid_234; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_749 = 8'heb == req_index | valid_235; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_750 = 8'hec == req_index | valid_236; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_751 = 8'hed == req_index | valid_237; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_752 = 8'hee == req_index | valid_238; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_753 = 8'hef == req_index | valid_239; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_754 = 8'hf0 == req_index | valid_240; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_755 = 8'hf1 == req_index | valid_241; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_756 = 8'hf2 == req_index | valid_242; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_757 = 8'hf3 == req_index | valid_243; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_758 = 8'hf4 == req_index | valid_244; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_759 = 8'hf5 == req_index | valid_245; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_760 = 8'hf6 == req_index | valid_246; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_761 = 8'hf7 == req_index | valid_247; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_762 = 8'hf8 == req_index | valid_248; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_763 = 8'hf9 == req_index | valid_249; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_764 = 8'hfa == req_index | valid_250; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_765 = 8'hfb == req_index | valid_251; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_766 = 8'hfc == req_index | valid_252; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_767 = 8'hfd == req_index | valid_253; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_768 = 8'hfe == req_index | valid_254; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire  _GEN_769 = 8'hff == req_index | valid_255; // @[Icache.scala 77:27 Icache.scala 77:27 Icache.scala 18:24]
  wire [19:0] _GEN_770 = 8'h0 == req_index ? req_tag : tag_0; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_771 = 8'h1 == req_index ? req_tag : tag_1; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_772 = 8'h2 == req_index ? req_tag : tag_2; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_773 = 8'h3 == req_index ? req_tag : tag_3; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_774 = 8'h4 == req_index ? req_tag : tag_4; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_775 = 8'h5 == req_index ? req_tag : tag_5; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_776 = 8'h6 == req_index ? req_tag : tag_6; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_777 = 8'h7 == req_index ? req_tag : tag_7; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_778 = 8'h8 == req_index ? req_tag : tag_8; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_779 = 8'h9 == req_index ? req_tag : tag_9; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_780 = 8'ha == req_index ? req_tag : tag_10; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_781 = 8'hb == req_index ? req_tag : tag_11; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_782 = 8'hc == req_index ? req_tag : tag_12; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_783 = 8'hd == req_index ? req_tag : tag_13; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_784 = 8'he == req_index ? req_tag : tag_14; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_785 = 8'hf == req_index ? req_tag : tag_15; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_786 = 8'h10 == req_index ? req_tag : tag_16; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_787 = 8'h11 == req_index ? req_tag : tag_17; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_788 = 8'h12 == req_index ? req_tag : tag_18; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_789 = 8'h13 == req_index ? req_tag : tag_19; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_790 = 8'h14 == req_index ? req_tag : tag_20; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_791 = 8'h15 == req_index ? req_tag : tag_21; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_792 = 8'h16 == req_index ? req_tag : tag_22; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_793 = 8'h17 == req_index ? req_tag : tag_23; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_794 = 8'h18 == req_index ? req_tag : tag_24; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_795 = 8'h19 == req_index ? req_tag : tag_25; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_796 = 8'h1a == req_index ? req_tag : tag_26; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_797 = 8'h1b == req_index ? req_tag : tag_27; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_798 = 8'h1c == req_index ? req_tag : tag_28; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_799 = 8'h1d == req_index ? req_tag : tag_29; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_800 = 8'h1e == req_index ? req_tag : tag_30; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_801 = 8'h1f == req_index ? req_tag : tag_31; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_802 = 8'h20 == req_index ? req_tag : tag_32; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_803 = 8'h21 == req_index ? req_tag : tag_33; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_804 = 8'h22 == req_index ? req_tag : tag_34; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_805 = 8'h23 == req_index ? req_tag : tag_35; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_806 = 8'h24 == req_index ? req_tag : tag_36; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_807 = 8'h25 == req_index ? req_tag : tag_37; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_808 = 8'h26 == req_index ? req_tag : tag_38; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_809 = 8'h27 == req_index ? req_tag : tag_39; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_810 = 8'h28 == req_index ? req_tag : tag_40; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_811 = 8'h29 == req_index ? req_tag : tag_41; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_812 = 8'h2a == req_index ? req_tag : tag_42; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_813 = 8'h2b == req_index ? req_tag : tag_43; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_814 = 8'h2c == req_index ? req_tag : tag_44; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_815 = 8'h2d == req_index ? req_tag : tag_45; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_816 = 8'h2e == req_index ? req_tag : tag_46; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_817 = 8'h2f == req_index ? req_tag : tag_47; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_818 = 8'h30 == req_index ? req_tag : tag_48; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_819 = 8'h31 == req_index ? req_tag : tag_49; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_820 = 8'h32 == req_index ? req_tag : tag_50; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_821 = 8'h33 == req_index ? req_tag : tag_51; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_822 = 8'h34 == req_index ? req_tag : tag_52; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_823 = 8'h35 == req_index ? req_tag : tag_53; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_824 = 8'h36 == req_index ? req_tag : tag_54; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_825 = 8'h37 == req_index ? req_tag : tag_55; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_826 = 8'h38 == req_index ? req_tag : tag_56; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_827 = 8'h39 == req_index ? req_tag : tag_57; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_828 = 8'h3a == req_index ? req_tag : tag_58; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_829 = 8'h3b == req_index ? req_tag : tag_59; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_830 = 8'h3c == req_index ? req_tag : tag_60; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_831 = 8'h3d == req_index ? req_tag : tag_61; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_832 = 8'h3e == req_index ? req_tag : tag_62; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_833 = 8'h3f == req_index ? req_tag : tag_63; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_834 = 8'h40 == req_index ? req_tag : tag_64; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_835 = 8'h41 == req_index ? req_tag : tag_65; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_836 = 8'h42 == req_index ? req_tag : tag_66; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_837 = 8'h43 == req_index ? req_tag : tag_67; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_838 = 8'h44 == req_index ? req_tag : tag_68; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_839 = 8'h45 == req_index ? req_tag : tag_69; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_840 = 8'h46 == req_index ? req_tag : tag_70; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_841 = 8'h47 == req_index ? req_tag : tag_71; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_842 = 8'h48 == req_index ? req_tag : tag_72; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_843 = 8'h49 == req_index ? req_tag : tag_73; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_844 = 8'h4a == req_index ? req_tag : tag_74; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_845 = 8'h4b == req_index ? req_tag : tag_75; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_846 = 8'h4c == req_index ? req_tag : tag_76; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_847 = 8'h4d == req_index ? req_tag : tag_77; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_848 = 8'h4e == req_index ? req_tag : tag_78; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_849 = 8'h4f == req_index ? req_tag : tag_79; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_850 = 8'h50 == req_index ? req_tag : tag_80; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_851 = 8'h51 == req_index ? req_tag : tag_81; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_852 = 8'h52 == req_index ? req_tag : tag_82; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_853 = 8'h53 == req_index ? req_tag : tag_83; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_854 = 8'h54 == req_index ? req_tag : tag_84; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_855 = 8'h55 == req_index ? req_tag : tag_85; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_856 = 8'h56 == req_index ? req_tag : tag_86; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_857 = 8'h57 == req_index ? req_tag : tag_87; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_858 = 8'h58 == req_index ? req_tag : tag_88; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_859 = 8'h59 == req_index ? req_tag : tag_89; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_860 = 8'h5a == req_index ? req_tag : tag_90; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_861 = 8'h5b == req_index ? req_tag : tag_91; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_862 = 8'h5c == req_index ? req_tag : tag_92; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_863 = 8'h5d == req_index ? req_tag : tag_93; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_864 = 8'h5e == req_index ? req_tag : tag_94; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_865 = 8'h5f == req_index ? req_tag : tag_95; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_866 = 8'h60 == req_index ? req_tag : tag_96; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_867 = 8'h61 == req_index ? req_tag : tag_97; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_868 = 8'h62 == req_index ? req_tag : tag_98; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_869 = 8'h63 == req_index ? req_tag : tag_99; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_870 = 8'h64 == req_index ? req_tag : tag_100; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_871 = 8'h65 == req_index ? req_tag : tag_101; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_872 = 8'h66 == req_index ? req_tag : tag_102; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_873 = 8'h67 == req_index ? req_tag : tag_103; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_874 = 8'h68 == req_index ? req_tag : tag_104; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_875 = 8'h69 == req_index ? req_tag : tag_105; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_876 = 8'h6a == req_index ? req_tag : tag_106; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_877 = 8'h6b == req_index ? req_tag : tag_107; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_878 = 8'h6c == req_index ? req_tag : tag_108; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_879 = 8'h6d == req_index ? req_tag : tag_109; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_880 = 8'h6e == req_index ? req_tag : tag_110; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_881 = 8'h6f == req_index ? req_tag : tag_111; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_882 = 8'h70 == req_index ? req_tag : tag_112; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_883 = 8'h71 == req_index ? req_tag : tag_113; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_884 = 8'h72 == req_index ? req_tag : tag_114; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_885 = 8'h73 == req_index ? req_tag : tag_115; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_886 = 8'h74 == req_index ? req_tag : tag_116; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_887 = 8'h75 == req_index ? req_tag : tag_117; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_888 = 8'h76 == req_index ? req_tag : tag_118; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_889 = 8'h77 == req_index ? req_tag : tag_119; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_890 = 8'h78 == req_index ? req_tag : tag_120; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_891 = 8'h79 == req_index ? req_tag : tag_121; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_892 = 8'h7a == req_index ? req_tag : tag_122; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_893 = 8'h7b == req_index ? req_tag : tag_123; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_894 = 8'h7c == req_index ? req_tag : tag_124; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_895 = 8'h7d == req_index ? req_tag : tag_125; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_896 = 8'h7e == req_index ? req_tag : tag_126; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_897 = 8'h7f == req_index ? req_tag : tag_127; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_898 = 8'h80 == req_index ? req_tag : tag_128; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_899 = 8'h81 == req_index ? req_tag : tag_129; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_900 = 8'h82 == req_index ? req_tag : tag_130; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_901 = 8'h83 == req_index ? req_tag : tag_131; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_902 = 8'h84 == req_index ? req_tag : tag_132; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_903 = 8'h85 == req_index ? req_tag : tag_133; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_904 = 8'h86 == req_index ? req_tag : tag_134; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_905 = 8'h87 == req_index ? req_tag : tag_135; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_906 = 8'h88 == req_index ? req_tag : tag_136; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_907 = 8'h89 == req_index ? req_tag : tag_137; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_908 = 8'h8a == req_index ? req_tag : tag_138; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_909 = 8'h8b == req_index ? req_tag : tag_139; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_910 = 8'h8c == req_index ? req_tag : tag_140; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_911 = 8'h8d == req_index ? req_tag : tag_141; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_912 = 8'h8e == req_index ? req_tag : tag_142; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_913 = 8'h8f == req_index ? req_tag : tag_143; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_914 = 8'h90 == req_index ? req_tag : tag_144; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_915 = 8'h91 == req_index ? req_tag : tag_145; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_916 = 8'h92 == req_index ? req_tag : tag_146; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_917 = 8'h93 == req_index ? req_tag : tag_147; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_918 = 8'h94 == req_index ? req_tag : tag_148; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_919 = 8'h95 == req_index ? req_tag : tag_149; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_920 = 8'h96 == req_index ? req_tag : tag_150; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_921 = 8'h97 == req_index ? req_tag : tag_151; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_922 = 8'h98 == req_index ? req_tag : tag_152; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_923 = 8'h99 == req_index ? req_tag : tag_153; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_924 = 8'h9a == req_index ? req_tag : tag_154; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_925 = 8'h9b == req_index ? req_tag : tag_155; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_926 = 8'h9c == req_index ? req_tag : tag_156; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_927 = 8'h9d == req_index ? req_tag : tag_157; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_928 = 8'h9e == req_index ? req_tag : tag_158; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_929 = 8'h9f == req_index ? req_tag : tag_159; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_930 = 8'ha0 == req_index ? req_tag : tag_160; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_931 = 8'ha1 == req_index ? req_tag : tag_161; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_932 = 8'ha2 == req_index ? req_tag : tag_162; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_933 = 8'ha3 == req_index ? req_tag : tag_163; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_934 = 8'ha4 == req_index ? req_tag : tag_164; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_935 = 8'ha5 == req_index ? req_tag : tag_165; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_936 = 8'ha6 == req_index ? req_tag : tag_166; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_937 = 8'ha7 == req_index ? req_tag : tag_167; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_938 = 8'ha8 == req_index ? req_tag : tag_168; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_939 = 8'ha9 == req_index ? req_tag : tag_169; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_940 = 8'haa == req_index ? req_tag : tag_170; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_941 = 8'hab == req_index ? req_tag : tag_171; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_942 = 8'hac == req_index ? req_tag : tag_172; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_943 = 8'had == req_index ? req_tag : tag_173; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_944 = 8'hae == req_index ? req_tag : tag_174; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_945 = 8'haf == req_index ? req_tag : tag_175; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_946 = 8'hb0 == req_index ? req_tag : tag_176; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_947 = 8'hb1 == req_index ? req_tag : tag_177; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_948 = 8'hb2 == req_index ? req_tag : tag_178; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_949 = 8'hb3 == req_index ? req_tag : tag_179; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_950 = 8'hb4 == req_index ? req_tag : tag_180; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_951 = 8'hb5 == req_index ? req_tag : tag_181; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_952 = 8'hb6 == req_index ? req_tag : tag_182; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_953 = 8'hb7 == req_index ? req_tag : tag_183; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_954 = 8'hb8 == req_index ? req_tag : tag_184; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_955 = 8'hb9 == req_index ? req_tag : tag_185; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_956 = 8'hba == req_index ? req_tag : tag_186; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_957 = 8'hbb == req_index ? req_tag : tag_187; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_958 = 8'hbc == req_index ? req_tag : tag_188; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_959 = 8'hbd == req_index ? req_tag : tag_189; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_960 = 8'hbe == req_index ? req_tag : tag_190; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_961 = 8'hbf == req_index ? req_tag : tag_191; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_962 = 8'hc0 == req_index ? req_tag : tag_192; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_963 = 8'hc1 == req_index ? req_tag : tag_193; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_964 = 8'hc2 == req_index ? req_tag : tag_194; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_965 = 8'hc3 == req_index ? req_tag : tag_195; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_966 = 8'hc4 == req_index ? req_tag : tag_196; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_967 = 8'hc5 == req_index ? req_tag : tag_197; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_968 = 8'hc6 == req_index ? req_tag : tag_198; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_969 = 8'hc7 == req_index ? req_tag : tag_199; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_970 = 8'hc8 == req_index ? req_tag : tag_200; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_971 = 8'hc9 == req_index ? req_tag : tag_201; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_972 = 8'hca == req_index ? req_tag : tag_202; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_973 = 8'hcb == req_index ? req_tag : tag_203; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_974 = 8'hcc == req_index ? req_tag : tag_204; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_975 = 8'hcd == req_index ? req_tag : tag_205; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_976 = 8'hce == req_index ? req_tag : tag_206; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_977 = 8'hcf == req_index ? req_tag : tag_207; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_978 = 8'hd0 == req_index ? req_tag : tag_208; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_979 = 8'hd1 == req_index ? req_tag : tag_209; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_980 = 8'hd2 == req_index ? req_tag : tag_210; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_981 = 8'hd3 == req_index ? req_tag : tag_211; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_982 = 8'hd4 == req_index ? req_tag : tag_212; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_983 = 8'hd5 == req_index ? req_tag : tag_213; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_984 = 8'hd6 == req_index ? req_tag : tag_214; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_985 = 8'hd7 == req_index ? req_tag : tag_215; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_986 = 8'hd8 == req_index ? req_tag : tag_216; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_987 = 8'hd9 == req_index ? req_tag : tag_217; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_988 = 8'hda == req_index ? req_tag : tag_218; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_989 = 8'hdb == req_index ? req_tag : tag_219; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_990 = 8'hdc == req_index ? req_tag : tag_220; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_991 = 8'hdd == req_index ? req_tag : tag_221; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_992 = 8'hde == req_index ? req_tag : tag_222; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_993 = 8'hdf == req_index ? req_tag : tag_223; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_994 = 8'he0 == req_index ? req_tag : tag_224; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_995 = 8'he1 == req_index ? req_tag : tag_225; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_996 = 8'he2 == req_index ? req_tag : tag_226; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_997 = 8'he3 == req_index ? req_tag : tag_227; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_998 = 8'he4 == req_index ? req_tag : tag_228; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_999 = 8'he5 == req_index ? req_tag : tag_229; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1000 = 8'he6 == req_index ? req_tag : tag_230; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1001 = 8'he7 == req_index ? req_tag : tag_231; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1002 = 8'he8 == req_index ? req_tag : tag_232; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1003 = 8'he9 == req_index ? req_tag : tag_233; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1004 = 8'hea == req_index ? req_tag : tag_234; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1005 = 8'heb == req_index ? req_tag : tag_235; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1006 = 8'hec == req_index ? req_tag : tag_236; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1007 = 8'hed == req_index ? req_tag : tag_237; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1008 = 8'hee == req_index ? req_tag : tag_238; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1009 = 8'hef == req_index ? req_tag : tag_239; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1010 = 8'hf0 == req_index ? req_tag : tag_240; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1011 = 8'hf1 == req_index ? req_tag : tag_241; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1012 = 8'hf2 == req_index ? req_tag : tag_242; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1013 = 8'hf3 == req_index ? req_tag : tag_243; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1014 = 8'hf4 == req_index ? req_tag : tag_244; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1015 = 8'hf5 == req_index ? req_tag : tag_245; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1016 = 8'hf6 == req_index ? req_tag : tag_246; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1017 = 8'hf7 == req_index ? req_tag : tag_247; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1018 = 8'hf8 == req_index ? req_tag : tag_248; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1019 = 8'hf9 == req_index ? req_tag : tag_249; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1020 = 8'hfa == req_index ? req_tag : tag_250; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1021 = 8'hfb == req_index ? req_tag : tag_251; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1022 = 8'hfc == req_index ? req_tag : tag_252; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1023 = 8'hfd == req_index ? req_tag : tag_253; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1024 = 8'hfe == req_index ? req_tag : tag_254; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire [19:0] _GEN_1025 = 8'hff == req_index ? req_tag : tag_255; // @[Icache.scala 78:27 Icache.scala 78:27 Icache.scala 17:24]
  wire  _GEN_1282 = cache_hit ? _GEN_514 : valid_0; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1283 = cache_hit ? _GEN_515 : valid_1; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1284 = cache_hit ? _GEN_516 : valid_2; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1285 = cache_hit ? _GEN_517 : valid_3; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1286 = cache_hit ? _GEN_518 : valid_4; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1287 = cache_hit ? _GEN_519 : valid_5; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1288 = cache_hit ? _GEN_520 : valid_6; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1289 = cache_hit ? _GEN_521 : valid_7; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1290 = cache_hit ? _GEN_522 : valid_8; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1291 = cache_hit ? _GEN_523 : valid_9; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1292 = cache_hit ? _GEN_524 : valid_10; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1293 = cache_hit ? _GEN_525 : valid_11; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1294 = cache_hit ? _GEN_526 : valid_12; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1295 = cache_hit ? _GEN_527 : valid_13; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1296 = cache_hit ? _GEN_528 : valid_14; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1297 = cache_hit ? _GEN_529 : valid_15; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1298 = cache_hit ? _GEN_530 : valid_16; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1299 = cache_hit ? _GEN_531 : valid_17; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1300 = cache_hit ? _GEN_532 : valid_18; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1301 = cache_hit ? _GEN_533 : valid_19; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1302 = cache_hit ? _GEN_534 : valid_20; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1303 = cache_hit ? _GEN_535 : valid_21; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1304 = cache_hit ? _GEN_536 : valid_22; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1305 = cache_hit ? _GEN_537 : valid_23; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1306 = cache_hit ? _GEN_538 : valid_24; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1307 = cache_hit ? _GEN_539 : valid_25; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1308 = cache_hit ? _GEN_540 : valid_26; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1309 = cache_hit ? _GEN_541 : valid_27; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1310 = cache_hit ? _GEN_542 : valid_28; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1311 = cache_hit ? _GEN_543 : valid_29; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1312 = cache_hit ? _GEN_544 : valid_30; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1313 = cache_hit ? _GEN_545 : valid_31; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1314 = cache_hit ? _GEN_546 : valid_32; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1315 = cache_hit ? _GEN_547 : valid_33; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1316 = cache_hit ? _GEN_548 : valid_34; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1317 = cache_hit ? _GEN_549 : valid_35; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1318 = cache_hit ? _GEN_550 : valid_36; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1319 = cache_hit ? _GEN_551 : valid_37; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1320 = cache_hit ? _GEN_552 : valid_38; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1321 = cache_hit ? _GEN_553 : valid_39; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1322 = cache_hit ? _GEN_554 : valid_40; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1323 = cache_hit ? _GEN_555 : valid_41; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1324 = cache_hit ? _GEN_556 : valid_42; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1325 = cache_hit ? _GEN_557 : valid_43; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1326 = cache_hit ? _GEN_558 : valid_44; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1327 = cache_hit ? _GEN_559 : valid_45; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1328 = cache_hit ? _GEN_560 : valid_46; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1329 = cache_hit ? _GEN_561 : valid_47; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1330 = cache_hit ? _GEN_562 : valid_48; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1331 = cache_hit ? _GEN_563 : valid_49; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1332 = cache_hit ? _GEN_564 : valid_50; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1333 = cache_hit ? _GEN_565 : valid_51; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1334 = cache_hit ? _GEN_566 : valid_52; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1335 = cache_hit ? _GEN_567 : valid_53; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1336 = cache_hit ? _GEN_568 : valid_54; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1337 = cache_hit ? _GEN_569 : valid_55; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1338 = cache_hit ? _GEN_570 : valid_56; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1339 = cache_hit ? _GEN_571 : valid_57; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1340 = cache_hit ? _GEN_572 : valid_58; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1341 = cache_hit ? _GEN_573 : valid_59; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1342 = cache_hit ? _GEN_574 : valid_60; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1343 = cache_hit ? _GEN_575 : valid_61; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1344 = cache_hit ? _GEN_576 : valid_62; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1345 = cache_hit ? _GEN_577 : valid_63; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1346 = cache_hit ? _GEN_578 : valid_64; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1347 = cache_hit ? _GEN_579 : valid_65; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1348 = cache_hit ? _GEN_580 : valid_66; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1349 = cache_hit ? _GEN_581 : valid_67; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1350 = cache_hit ? _GEN_582 : valid_68; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1351 = cache_hit ? _GEN_583 : valid_69; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1352 = cache_hit ? _GEN_584 : valid_70; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1353 = cache_hit ? _GEN_585 : valid_71; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1354 = cache_hit ? _GEN_586 : valid_72; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1355 = cache_hit ? _GEN_587 : valid_73; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1356 = cache_hit ? _GEN_588 : valid_74; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1357 = cache_hit ? _GEN_589 : valid_75; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1358 = cache_hit ? _GEN_590 : valid_76; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1359 = cache_hit ? _GEN_591 : valid_77; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1360 = cache_hit ? _GEN_592 : valid_78; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1361 = cache_hit ? _GEN_593 : valid_79; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1362 = cache_hit ? _GEN_594 : valid_80; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1363 = cache_hit ? _GEN_595 : valid_81; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1364 = cache_hit ? _GEN_596 : valid_82; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1365 = cache_hit ? _GEN_597 : valid_83; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1366 = cache_hit ? _GEN_598 : valid_84; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1367 = cache_hit ? _GEN_599 : valid_85; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1368 = cache_hit ? _GEN_600 : valid_86; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1369 = cache_hit ? _GEN_601 : valid_87; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1370 = cache_hit ? _GEN_602 : valid_88; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1371 = cache_hit ? _GEN_603 : valid_89; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1372 = cache_hit ? _GEN_604 : valid_90; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1373 = cache_hit ? _GEN_605 : valid_91; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1374 = cache_hit ? _GEN_606 : valid_92; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1375 = cache_hit ? _GEN_607 : valid_93; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1376 = cache_hit ? _GEN_608 : valid_94; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1377 = cache_hit ? _GEN_609 : valid_95; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1378 = cache_hit ? _GEN_610 : valid_96; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1379 = cache_hit ? _GEN_611 : valid_97; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1380 = cache_hit ? _GEN_612 : valid_98; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1381 = cache_hit ? _GEN_613 : valid_99; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1382 = cache_hit ? _GEN_614 : valid_100; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1383 = cache_hit ? _GEN_615 : valid_101; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1384 = cache_hit ? _GEN_616 : valid_102; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1385 = cache_hit ? _GEN_617 : valid_103; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1386 = cache_hit ? _GEN_618 : valid_104; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1387 = cache_hit ? _GEN_619 : valid_105; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1388 = cache_hit ? _GEN_620 : valid_106; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1389 = cache_hit ? _GEN_621 : valid_107; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1390 = cache_hit ? _GEN_622 : valid_108; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1391 = cache_hit ? _GEN_623 : valid_109; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1392 = cache_hit ? _GEN_624 : valid_110; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1393 = cache_hit ? _GEN_625 : valid_111; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1394 = cache_hit ? _GEN_626 : valid_112; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1395 = cache_hit ? _GEN_627 : valid_113; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1396 = cache_hit ? _GEN_628 : valid_114; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1397 = cache_hit ? _GEN_629 : valid_115; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1398 = cache_hit ? _GEN_630 : valid_116; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1399 = cache_hit ? _GEN_631 : valid_117; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1400 = cache_hit ? _GEN_632 : valid_118; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1401 = cache_hit ? _GEN_633 : valid_119; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1402 = cache_hit ? _GEN_634 : valid_120; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1403 = cache_hit ? _GEN_635 : valid_121; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1404 = cache_hit ? _GEN_636 : valid_122; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1405 = cache_hit ? _GEN_637 : valid_123; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1406 = cache_hit ? _GEN_638 : valid_124; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1407 = cache_hit ? _GEN_639 : valid_125; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1408 = cache_hit ? _GEN_640 : valid_126; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1409 = cache_hit ? _GEN_641 : valid_127; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1410 = cache_hit ? _GEN_642 : valid_128; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1411 = cache_hit ? _GEN_643 : valid_129; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1412 = cache_hit ? _GEN_644 : valid_130; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1413 = cache_hit ? _GEN_645 : valid_131; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1414 = cache_hit ? _GEN_646 : valid_132; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1415 = cache_hit ? _GEN_647 : valid_133; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1416 = cache_hit ? _GEN_648 : valid_134; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1417 = cache_hit ? _GEN_649 : valid_135; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1418 = cache_hit ? _GEN_650 : valid_136; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1419 = cache_hit ? _GEN_651 : valid_137; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1420 = cache_hit ? _GEN_652 : valid_138; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1421 = cache_hit ? _GEN_653 : valid_139; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1422 = cache_hit ? _GEN_654 : valid_140; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1423 = cache_hit ? _GEN_655 : valid_141; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1424 = cache_hit ? _GEN_656 : valid_142; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1425 = cache_hit ? _GEN_657 : valid_143; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1426 = cache_hit ? _GEN_658 : valid_144; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1427 = cache_hit ? _GEN_659 : valid_145; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1428 = cache_hit ? _GEN_660 : valid_146; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1429 = cache_hit ? _GEN_661 : valid_147; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1430 = cache_hit ? _GEN_662 : valid_148; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1431 = cache_hit ? _GEN_663 : valid_149; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1432 = cache_hit ? _GEN_664 : valid_150; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1433 = cache_hit ? _GEN_665 : valid_151; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1434 = cache_hit ? _GEN_666 : valid_152; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1435 = cache_hit ? _GEN_667 : valid_153; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1436 = cache_hit ? _GEN_668 : valid_154; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1437 = cache_hit ? _GEN_669 : valid_155; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1438 = cache_hit ? _GEN_670 : valid_156; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1439 = cache_hit ? _GEN_671 : valid_157; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1440 = cache_hit ? _GEN_672 : valid_158; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1441 = cache_hit ? _GEN_673 : valid_159; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1442 = cache_hit ? _GEN_674 : valid_160; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1443 = cache_hit ? _GEN_675 : valid_161; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1444 = cache_hit ? _GEN_676 : valid_162; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1445 = cache_hit ? _GEN_677 : valid_163; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1446 = cache_hit ? _GEN_678 : valid_164; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1447 = cache_hit ? _GEN_679 : valid_165; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1448 = cache_hit ? _GEN_680 : valid_166; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1449 = cache_hit ? _GEN_681 : valid_167; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1450 = cache_hit ? _GEN_682 : valid_168; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1451 = cache_hit ? _GEN_683 : valid_169; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1452 = cache_hit ? _GEN_684 : valid_170; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1453 = cache_hit ? _GEN_685 : valid_171; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1454 = cache_hit ? _GEN_686 : valid_172; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1455 = cache_hit ? _GEN_687 : valid_173; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1456 = cache_hit ? _GEN_688 : valid_174; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1457 = cache_hit ? _GEN_689 : valid_175; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1458 = cache_hit ? _GEN_690 : valid_176; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1459 = cache_hit ? _GEN_691 : valid_177; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1460 = cache_hit ? _GEN_692 : valid_178; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1461 = cache_hit ? _GEN_693 : valid_179; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1462 = cache_hit ? _GEN_694 : valid_180; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1463 = cache_hit ? _GEN_695 : valid_181; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1464 = cache_hit ? _GEN_696 : valid_182; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1465 = cache_hit ? _GEN_697 : valid_183; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1466 = cache_hit ? _GEN_698 : valid_184; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1467 = cache_hit ? _GEN_699 : valid_185; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1468 = cache_hit ? _GEN_700 : valid_186; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1469 = cache_hit ? _GEN_701 : valid_187; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1470 = cache_hit ? _GEN_702 : valid_188; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1471 = cache_hit ? _GEN_703 : valid_189; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1472 = cache_hit ? _GEN_704 : valid_190; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1473 = cache_hit ? _GEN_705 : valid_191; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1474 = cache_hit ? _GEN_706 : valid_192; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1475 = cache_hit ? _GEN_707 : valid_193; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1476 = cache_hit ? _GEN_708 : valid_194; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1477 = cache_hit ? _GEN_709 : valid_195; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1478 = cache_hit ? _GEN_710 : valid_196; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1479 = cache_hit ? _GEN_711 : valid_197; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1480 = cache_hit ? _GEN_712 : valid_198; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1481 = cache_hit ? _GEN_713 : valid_199; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1482 = cache_hit ? _GEN_714 : valid_200; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1483 = cache_hit ? _GEN_715 : valid_201; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1484 = cache_hit ? _GEN_716 : valid_202; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1485 = cache_hit ? _GEN_717 : valid_203; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1486 = cache_hit ? _GEN_718 : valid_204; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1487 = cache_hit ? _GEN_719 : valid_205; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1488 = cache_hit ? _GEN_720 : valid_206; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1489 = cache_hit ? _GEN_721 : valid_207; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1490 = cache_hit ? _GEN_722 : valid_208; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1491 = cache_hit ? _GEN_723 : valid_209; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1492 = cache_hit ? _GEN_724 : valid_210; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1493 = cache_hit ? _GEN_725 : valid_211; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1494 = cache_hit ? _GEN_726 : valid_212; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1495 = cache_hit ? _GEN_727 : valid_213; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1496 = cache_hit ? _GEN_728 : valid_214; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1497 = cache_hit ? _GEN_729 : valid_215; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1498 = cache_hit ? _GEN_730 : valid_216; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1499 = cache_hit ? _GEN_731 : valid_217; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1500 = cache_hit ? _GEN_732 : valid_218; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1501 = cache_hit ? _GEN_733 : valid_219; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1502 = cache_hit ? _GEN_734 : valid_220; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1503 = cache_hit ? _GEN_735 : valid_221; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1504 = cache_hit ? _GEN_736 : valid_222; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1505 = cache_hit ? _GEN_737 : valid_223; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1506 = cache_hit ? _GEN_738 : valid_224; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1507 = cache_hit ? _GEN_739 : valid_225; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1508 = cache_hit ? _GEN_740 : valid_226; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1509 = cache_hit ? _GEN_741 : valid_227; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1510 = cache_hit ? _GEN_742 : valid_228; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1511 = cache_hit ? _GEN_743 : valid_229; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1512 = cache_hit ? _GEN_744 : valid_230; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1513 = cache_hit ? _GEN_745 : valid_231; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1514 = cache_hit ? _GEN_746 : valid_232; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1515 = cache_hit ? _GEN_747 : valid_233; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1516 = cache_hit ? _GEN_748 : valid_234; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1517 = cache_hit ? _GEN_749 : valid_235; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1518 = cache_hit ? _GEN_750 : valid_236; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1519 = cache_hit ? _GEN_751 : valid_237; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1520 = cache_hit ? _GEN_752 : valid_238; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1521 = cache_hit ? _GEN_753 : valid_239; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1522 = cache_hit ? _GEN_754 : valid_240; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1523 = cache_hit ? _GEN_755 : valid_241; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1524 = cache_hit ? _GEN_756 : valid_242; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1525 = cache_hit ? _GEN_757 : valid_243; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1526 = cache_hit ? _GEN_758 : valid_244; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1527 = cache_hit ? _GEN_759 : valid_245; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1528 = cache_hit ? _GEN_760 : valid_246; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1529 = cache_hit ? _GEN_761 : valid_247; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1530 = cache_hit ? _GEN_762 : valid_248; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1531 = cache_hit ? _GEN_763 : valid_249; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1532 = cache_hit ? _GEN_764 : valid_250; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1533 = cache_hit ? _GEN_765 : valid_251; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1534 = cache_hit ? _GEN_766 : valid_252; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1535 = cache_hit ? _GEN_767 : valid_253; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1536 = cache_hit ? _GEN_768 : valid_254; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire  _GEN_1537 = cache_hit ? _GEN_769 : valid_255; // @[Icache.scala 76:29 Icache.scala 18:24]
  wire [19:0] _GEN_1538 = cache_hit ? _GEN_770 : tag_0; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1539 = cache_hit ? _GEN_771 : tag_1; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1540 = cache_hit ? _GEN_772 : tag_2; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1541 = cache_hit ? _GEN_773 : tag_3; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1542 = cache_hit ? _GEN_774 : tag_4; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1543 = cache_hit ? _GEN_775 : tag_5; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1544 = cache_hit ? _GEN_776 : tag_6; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1545 = cache_hit ? _GEN_777 : tag_7; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1546 = cache_hit ? _GEN_778 : tag_8; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1547 = cache_hit ? _GEN_779 : tag_9; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1548 = cache_hit ? _GEN_780 : tag_10; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1549 = cache_hit ? _GEN_781 : tag_11; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1550 = cache_hit ? _GEN_782 : tag_12; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1551 = cache_hit ? _GEN_783 : tag_13; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1552 = cache_hit ? _GEN_784 : tag_14; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1553 = cache_hit ? _GEN_785 : tag_15; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1554 = cache_hit ? _GEN_786 : tag_16; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1555 = cache_hit ? _GEN_787 : tag_17; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1556 = cache_hit ? _GEN_788 : tag_18; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1557 = cache_hit ? _GEN_789 : tag_19; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1558 = cache_hit ? _GEN_790 : tag_20; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1559 = cache_hit ? _GEN_791 : tag_21; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1560 = cache_hit ? _GEN_792 : tag_22; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1561 = cache_hit ? _GEN_793 : tag_23; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1562 = cache_hit ? _GEN_794 : tag_24; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1563 = cache_hit ? _GEN_795 : tag_25; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1564 = cache_hit ? _GEN_796 : tag_26; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1565 = cache_hit ? _GEN_797 : tag_27; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1566 = cache_hit ? _GEN_798 : tag_28; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1567 = cache_hit ? _GEN_799 : tag_29; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1568 = cache_hit ? _GEN_800 : tag_30; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1569 = cache_hit ? _GEN_801 : tag_31; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1570 = cache_hit ? _GEN_802 : tag_32; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1571 = cache_hit ? _GEN_803 : tag_33; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1572 = cache_hit ? _GEN_804 : tag_34; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1573 = cache_hit ? _GEN_805 : tag_35; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1574 = cache_hit ? _GEN_806 : tag_36; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1575 = cache_hit ? _GEN_807 : tag_37; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1576 = cache_hit ? _GEN_808 : tag_38; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1577 = cache_hit ? _GEN_809 : tag_39; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1578 = cache_hit ? _GEN_810 : tag_40; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1579 = cache_hit ? _GEN_811 : tag_41; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1580 = cache_hit ? _GEN_812 : tag_42; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1581 = cache_hit ? _GEN_813 : tag_43; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1582 = cache_hit ? _GEN_814 : tag_44; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1583 = cache_hit ? _GEN_815 : tag_45; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1584 = cache_hit ? _GEN_816 : tag_46; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1585 = cache_hit ? _GEN_817 : tag_47; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1586 = cache_hit ? _GEN_818 : tag_48; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1587 = cache_hit ? _GEN_819 : tag_49; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1588 = cache_hit ? _GEN_820 : tag_50; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1589 = cache_hit ? _GEN_821 : tag_51; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1590 = cache_hit ? _GEN_822 : tag_52; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1591 = cache_hit ? _GEN_823 : tag_53; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1592 = cache_hit ? _GEN_824 : tag_54; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1593 = cache_hit ? _GEN_825 : tag_55; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1594 = cache_hit ? _GEN_826 : tag_56; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1595 = cache_hit ? _GEN_827 : tag_57; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1596 = cache_hit ? _GEN_828 : tag_58; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1597 = cache_hit ? _GEN_829 : tag_59; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1598 = cache_hit ? _GEN_830 : tag_60; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1599 = cache_hit ? _GEN_831 : tag_61; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1600 = cache_hit ? _GEN_832 : tag_62; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1601 = cache_hit ? _GEN_833 : tag_63; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1602 = cache_hit ? _GEN_834 : tag_64; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1603 = cache_hit ? _GEN_835 : tag_65; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1604 = cache_hit ? _GEN_836 : tag_66; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1605 = cache_hit ? _GEN_837 : tag_67; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1606 = cache_hit ? _GEN_838 : tag_68; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1607 = cache_hit ? _GEN_839 : tag_69; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1608 = cache_hit ? _GEN_840 : tag_70; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1609 = cache_hit ? _GEN_841 : tag_71; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1610 = cache_hit ? _GEN_842 : tag_72; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1611 = cache_hit ? _GEN_843 : tag_73; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1612 = cache_hit ? _GEN_844 : tag_74; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1613 = cache_hit ? _GEN_845 : tag_75; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1614 = cache_hit ? _GEN_846 : tag_76; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1615 = cache_hit ? _GEN_847 : tag_77; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1616 = cache_hit ? _GEN_848 : tag_78; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1617 = cache_hit ? _GEN_849 : tag_79; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1618 = cache_hit ? _GEN_850 : tag_80; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1619 = cache_hit ? _GEN_851 : tag_81; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1620 = cache_hit ? _GEN_852 : tag_82; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1621 = cache_hit ? _GEN_853 : tag_83; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1622 = cache_hit ? _GEN_854 : tag_84; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1623 = cache_hit ? _GEN_855 : tag_85; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1624 = cache_hit ? _GEN_856 : tag_86; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1625 = cache_hit ? _GEN_857 : tag_87; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1626 = cache_hit ? _GEN_858 : tag_88; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1627 = cache_hit ? _GEN_859 : tag_89; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1628 = cache_hit ? _GEN_860 : tag_90; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1629 = cache_hit ? _GEN_861 : tag_91; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1630 = cache_hit ? _GEN_862 : tag_92; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1631 = cache_hit ? _GEN_863 : tag_93; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1632 = cache_hit ? _GEN_864 : tag_94; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1633 = cache_hit ? _GEN_865 : tag_95; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1634 = cache_hit ? _GEN_866 : tag_96; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1635 = cache_hit ? _GEN_867 : tag_97; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1636 = cache_hit ? _GEN_868 : tag_98; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1637 = cache_hit ? _GEN_869 : tag_99; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1638 = cache_hit ? _GEN_870 : tag_100; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1639 = cache_hit ? _GEN_871 : tag_101; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1640 = cache_hit ? _GEN_872 : tag_102; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1641 = cache_hit ? _GEN_873 : tag_103; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1642 = cache_hit ? _GEN_874 : tag_104; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1643 = cache_hit ? _GEN_875 : tag_105; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1644 = cache_hit ? _GEN_876 : tag_106; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1645 = cache_hit ? _GEN_877 : tag_107; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1646 = cache_hit ? _GEN_878 : tag_108; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1647 = cache_hit ? _GEN_879 : tag_109; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1648 = cache_hit ? _GEN_880 : tag_110; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1649 = cache_hit ? _GEN_881 : tag_111; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1650 = cache_hit ? _GEN_882 : tag_112; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1651 = cache_hit ? _GEN_883 : tag_113; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1652 = cache_hit ? _GEN_884 : tag_114; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1653 = cache_hit ? _GEN_885 : tag_115; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1654 = cache_hit ? _GEN_886 : tag_116; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1655 = cache_hit ? _GEN_887 : tag_117; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1656 = cache_hit ? _GEN_888 : tag_118; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1657 = cache_hit ? _GEN_889 : tag_119; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1658 = cache_hit ? _GEN_890 : tag_120; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1659 = cache_hit ? _GEN_891 : tag_121; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1660 = cache_hit ? _GEN_892 : tag_122; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1661 = cache_hit ? _GEN_893 : tag_123; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1662 = cache_hit ? _GEN_894 : tag_124; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1663 = cache_hit ? _GEN_895 : tag_125; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1664 = cache_hit ? _GEN_896 : tag_126; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1665 = cache_hit ? _GEN_897 : tag_127; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1666 = cache_hit ? _GEN_898 : tag_128; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1667 = cache_hit ? _GEN_899 : tag_129; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1668 = cache_hit ? _GEN_900 : tag_130; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1669 = cache_hit ? _GEN_901 : tag_131; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1670 = cache_hit ? _GEN_902 : tag_132; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1671 = cache_hit ? _GEN_903 : tag_133; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1672 = cache_hit ? _GEN_904 : tag_134; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1673 = cache_hit ? _GEN_905 : tag_135; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1674 = cache_hit ? _GEN_906 : tag_136; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1675 = cache_hit ? _GEN_907 : tag_137; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1676 = cache_hit ? _GEN_908 : tag_138; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1677 = cache_hit ? _GEN_909 : tag_139; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1678 = cache_hit ? _GEN_910 : tag_140; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1679 = cache_hit ? _GEN_911 : tag_141; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1680 = cache_hit ? _GEN_912 : tag_142; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1681 = cache_hit ? _GEN_913 : tag_143; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1682 = cache_hit ? _GEN_914 : tag_144; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1683 = cache_hit ? _GEN_915 : tag_145; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1684 = cache_hit ? _GEN_916 : tag_146; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1685 = cache_hit ? _GEN_917 : tag_147; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1686 = cache_hit ? _GEN_918 : tag_148; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1687 = cache_hit ? _GEN_919 : tag_149; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1688 = cache_hit ? _GEN_920 : tag_150; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1689 = cache_hit ? _GEN_921 : tag_151; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1690 = cache_hit ? _GEN_922 : tag_152; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1691 = cache_hit ? _GEN_923 : tag_153; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1692 = cache_hit ? _GEN_924 : tag_154; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1693 = cache_hit ? _GEN_925 : tag_155; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1694 = cache_hit ? _GEN_926 : tag_156; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1695 = cache_hit ? _GEN_927 : tag_157; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1696 = cache_hit ? _GEN_928 : tag_158; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1697 = cache_hit ? _GEN_929 : tag_159; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1698 = cache_hit ? _GEN_930 : tag_160; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1699 = cache_hit ? _GEN_931 : tag_161; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1700 = cache_hit ? _GEN_932 : tag_162; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1701 = cache_hit ? _GEN_933 : tag_163; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1702 = cache_hit ? _GEN_934 : tag_164; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1703 = cache_hit ? _GEN_935 : tag_165; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1704 = cache_hit ? _GEN_936 : tag_166; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1705 = cache_hit ? _GEN_937 : tag_167; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1706 = cache_hit ? _GEN_938 : tag_168; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1707 = cache_hit ? _GEN_939 : tag_169; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1708 = cache_hit ? _GEN_940 : tag_170; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1709 = cache_hit ? _GEN_941 : tag_171; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1710 = cache_hit ? _GEN_942 : tag_172; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1711 = cache_hit ? _GEN_943 : tag_173; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1712 = cache_hit ? _GEN_944 : tag_174; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1713 = cache_hit ? _GEN_945 : tag_175; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1714 = cache_hit ? _GEN_946 : tag_176; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1715 = cache_hit ? _GEN_947 : tag_177; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1716 = cache_hit ? _GEN_948 : tag_178; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1717 = cache_hit ? _GEN_949 : tag_179; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1718 = cache_hit ? _GEN_950 : tag_180; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1719 = cache_hit ? _GEN_951 : tag_181; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1720 = cache_hit ? _GEN_952 : tag_182; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1721 = cache_hit ? _GEN_953 : tag_183; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1722 = cache_hit ? _GEN_954 : tag_184; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1723 = cache_hit ? _GEN_955 : tag_185; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1724 = cache_hit ? _GEN_956 : tag_186; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1725 = cache_hit ? _GEN_957 : tag_187; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1726 = cache_hit ? _GEN_958 : tag_188; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1727 = cache_hit ? _GEN_959 : tag_189; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1728 = cache_hit ? _GEN_960 : tag_190; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1729 = cache_hit ? _GEN_961 : tag_191; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1730 = cache_hit ? _GEN_962 : tag_192; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1731 = cache_hit ? _GEN_963 : tag_193; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1732 = cache_hit ? _GEN_964 : tag_194; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1733 = cache_hit ? _GEN_965 : tag_195; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1734 = cache_hit ? _GEN_966 : tag_196; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1735 = cache_hit ? _GEN_967 : tag_197; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1736 = cache_hit ? _GEN_968 : tag_198; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1737 = cache_hit ? _GEN_969 : tag_199; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1738 = cache_hit ? _GEN_970 : tag_200; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1739 = cache_hit ? _GEN_971 : tag_201; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1740 = cache_hit ? _GEN_972 : tag_202; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1741 = cache_hit ? _GEN_973 : tag_203; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1742 = cache_hit ? _GEN_974 : tag_204; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1743 = cache_hit ? _GEN_975 : tag_205; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1744 = cache_hit ? _GEN_976 : tag_206; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1745 = cache_hit ? _GEN_977 : tag_207; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1746 = cache_hit ? _GEN_978 : tag_208; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1747 = cache_hit ? _GEN_979 : tag_209; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1748 = cache_hit ? _GEN_980 : tag_210; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1749 = cache_hit ? _GEN_981 : tag_211; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1750 = cache_hit ? _GEN_982 : tag_212; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1751 = cache_hit ? _GEN_983 : tag_213; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1752 = cache_hit ? _GEN_984 : tag_214; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1753 = cache_hit ? _GEN_985 : tag_215; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1754 = cache_hit ? _GEN_986 : tag_216; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1755 = cache_hit ? _GEN_987 : tag_217; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1756 = cache_hit ? _GEN_988 : tag_218; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1757 = cache_hit ? _GEN_989 : tag_219; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1758 = cache_hit ? _GEN_990 : tag_220; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1759 = cache_hit ? _GEN_991 : tag_221; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1760 = cache_hit ? _GEN_992 : tag_222; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1761 = cache_hit ? _GEN_993 : tag_223; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1762 = cache_hit ? _GEN_994 : tag_224; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1763 = cache_hit ? _GEN_995 : tag_225; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1764 = cache_hit ? _GEN_996 : tag_226; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1765 = cache_hit ? _GEN_997 : tag_227; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1766 = cache_hit ? _GEN_998 : tag_228; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1767 = cache_hit ? _GEN_999 : tag_229; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1768 = cache_hit ? _GEN_1000 : tag_230; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1769 = cache_hit ? _GEN_1001 : tag_231; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1770 = cache_hit ? _GEN_1002 : tag_232; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1771 = cache_hit ? _GEN_1003 : tag_233; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1772 = cache_hit ? _GEN_1004 : tag_234; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1773 = cache_hit ? _GEN_1005 : tag_235; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1774 = cache_hit ? _GEN_1006 : tag_236; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1775 = cache_hit ? _GEN_1007 : tag_237; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1776 = cache_hit ? _GEN_1008 : tag_238; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1777 = cache_hit ? _GEN_1009 : tag_239; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1778 = cache_hit ? _GEN_1010 : tag_240; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1779 = cache_hit ? _GEN_1011 : tag_241; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1780 = cache_hit ? _GEN_1012 : tag_242; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1781 = cache_hit ? _GEN_1013 : tag_243; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1782 = cache_hit ? _GEN_1014 : tag_244; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1783 = cache_hit ? _GEN_1015 : tag_245; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1784 = cache_hit ? _GEN_1016 : tag_246; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1785 = cache_hit ? _GEN_1017 : tag_247; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1786 = cache_hit ? _GEN_1018 : tag_248; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1787 = cache_hit ? _GEN_1019 : tag_249; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1788 = cache_hit ? _GEN_1020 : tag_250; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1789 = cache_hit ? _GEN_1021 : tag_251; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1790 = cache_hit ? _GEN_1022 : tag_252; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1791 = cache_hit ? _GEN_1023 : tag_253; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1792 = cache_hit ? _GEN_1024 : tag_254; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire [19:0] _GEN_1793 = cache_hit ? _GEN_1025 : tag_255; // @[Icache.scala 76:29 Icache.scala 17:24]
  wire  _GEN_2050 = cache_hit | inst_ready; // @[Icache.scala 76:29 Icache.scala 80:27 Icache.scala 42:28]
  wire [2:0] _GEN_2051 = cache_hit ? 3'h0 : 3'h3; // @[Icache.scala 76:29 Icache.scala 81:27 Icache.scala 84:21]
  wire [2:0] _GEN_2052 = io_br_stall ? 3'h0 : _GEN_2051; // @[Icache.scala 73:26 Icache.scala 74:15]
  wire  _GEN_2053 = io_br_stall ? valid_0 : _GEN_1282; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2054 = io_br_stall ? valid_1 : _GEN_1283; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2055 = io_br_stall ? valid_2 : _GEN_1284; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2056 = io_br_stall ? valid_3 : _GEN_1285; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2057 = io_br_stall ? valid_4 : _GEN_1286; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2058 = io_br_stall ? valid_5 : _GEN_1287; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2059 = io_br_stall ? valid_6 : _GEN_1288; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2060 = io_br_stall ? valid_7 : _GEN_1289; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2061 = io_br_stall ? valid_8 : _GEN_1290; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2062 = io_br_stall ? valid_9 : _GEN_1291; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2063 = io_br_stall ? valid_10 : _GEN_1292; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2064 = io_br_stall ? valid_11 : _GEN_1293; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2065 = io_br_stall ? valid_12 : _GEN_1294; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2066 = io_br_stall ? valid_13 : _GEN_1295; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2067 = io_br_stall ? valid_14 : _GEN_1296; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2068 = io_br_stall ? valid_15 : _GEN_1297; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2069 = io_br_stall ? valid_16 : _GEN_1298; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2070 = io_br_stall ? valid_17 : _GEN_1299; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2071 = io_br_stall ? valid_18 : _GEN_1300; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2072 = io_br_stall ? valid_19 : _GEN_1301; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2073 = io_br_stall ? valid_20 : _GEN_1302; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2074 = io_br_stall ? valid_21 : _GEN_1303; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2075 = io_br_stall ? valid_22 : _GEN_1304; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2076 = io_br_stall ? valid_23 : _GEN_1305; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2077 = io_br_stall ? valid_24 : _GEN_1306; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2078 = io_br_stall ? valid_25 : _GEN_1307; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2079 = io_br_stall ? valid_26 : _GEN_1308; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2080 = io_br_stall ? valid_27 : _GEN_1309; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2081 = io_br_stall ? valid_28 : _GEN_1310; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2082 = io_br_stall ? valid_29 : _GEN_1311; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2083 = io_br_stall ? valid_30 : _GEN_1312; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2084 = io_br_stall ? valid_31 : _GEN_1313; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2085 = io_br_stall ? valid_32 : _GEN_1314; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2086 = io_br_stall ? valid_33 : _GEN_1315; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2087 = io_br_stall ? valid_34 : _GEN_1316; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2088 = io_br_stall ? valid_35 : _GEN_1317; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2089 = io_br_stall ? valid_36 : _GEN_1318; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2090 = io_br_stall ? valid_37 : _GEN_1319; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2091 = io_br_stall ? valid_38 : _GEN_1320; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2092 = io_br_stall ? valid_39 : _GEN_1321; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2093 = io_br_stall ? valid_40 : _GEN_1322; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2094 = io_br_stall ? valid_41 : _GEN_1323; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2095 = io_br_stall ? valid_42 : _GEN_1324; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2096 = io_br_stall ? valid_43 : _GEN_1325; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2097 = io_br_stall ? valid_44 : _GEN_1326; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2098 = io_br_stall ? valid_45 : _GEN_1327; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2099 = io_br_stall ? valid_46 : _GEN_1328; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2100 = io_br_stall ? valid_47 : _GEN_1329; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2101 = io_br_stall ? valid_48 : _GEN_1330; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2102 = io_br_stall ? valid_49 : _GEN_1331; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2103 = io_br_stall ? valid_50 : _GEN_1332; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2104 = io_br_stall ? valid_51 : _GEN_1333; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2105 = io_br_stall ? valid_52 : _GEN_1334; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2106 = io_br_stall ? valid_53 : _GEN_1335; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2107 = io_br_stall ? valid_54 : _GEN_1336; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2108 = io_br_stall ? valid_55 : _GEN_1337; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2109 = io_br_stall ? valid_56 : _GEN_1338; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2110 = io_br_stall ? valid_57 : _GEN_1339; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2111 = io_br_stall ? valid_58 : _GEN_1340; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2112 = io_br_stall ? valid_59 : _GEN_1341; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2113 = io_br_stall ? valid_60 : _GEN_1342; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2114 = io_br_stall ? valid_61 : _GEN_1343; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2115 = io_br_stall ? valid_62 : _GEN_1344; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2116 = io_br_stall ? valid_63 : _GEN_1345; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2117 = io_br_stall ? valid_64 : _GEN_1346; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2118 = io_br_stall ? valid_65 : _GEN_1347; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2119 = io_br_stall ? valid_66 : _GEN_1348; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2120 = io_br_stall ? valid_67 : _GEN_1349; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2121 = io_br_stall ? valid_68 : _GEN_1350; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2122 = io_br_stall ? valid_69 : _GEN_1351; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2123 = io_br_stall ? valid_70 : _GEN_1352; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2124 = io_br_stall ? valid_71 : _GEN_1353; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2125 = io_br_stall ? valid_72 : _GEN_1354; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2126 = io_br_stall ? valid_73 : _GEN_1355; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2127 = io_br_stall ? valid_74 : _GEN_1356; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2128 = io_br_stall ? valid_75 : _GEN_1357; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2129 = io_br_stall ? valid_76 : _GEN_1358; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2130 = io_br_stall ? valid_77 : _GEN_1359; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2131 = io_br_stall ? valid_78 : _GEN_1360; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2132 = io_br_stall ? valid_79 : _GEN_1361; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2133 = io_br_stall ? valid_80 : _GEN_1362; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2134 = io_br_stall ? valid_81 : _GEN_1363; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2135 = io_br_stall ? valid_82 : _GEN_1364; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2136 = io_br_stall ? valid_83 : _GEN_1365; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2137 = io_br_stall ? valid_84 : _GEN_1366; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2138 = io_br_stall ? valid_85 : _GEN_1367; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2139 = io_br_stall ? valid_86 : _GEN_1368; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2140 = io_br_stall ? valid_87 : _GEN_1369; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2141 = io_br_stall ? valid_88 : _GEN_1370; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2142 = io_br_stall ? valid_89 : _GEN_1371; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2143 = io_br_stall ? valid_90 : _GEN_1372; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2144 = io_br_stall ? valid_91 : _GEN_1373; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2145 = io_br_stall ? valid_92 : _GEN_1374; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2146 = io_br_stall ? valid_93 : _GEN_1375; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2147 = io_br_stall ? valid_94 : _GEN_1376; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2148 = io_br_stall ? valid_95 : _GEN_1377; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2149 = io_br_stall ? valid_96 : _GEN_1378; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2150 = io_br_stall ? valid_97 : _GEN_1379; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2151 = io_br_stall ? valid_98 : _GEN_1380; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2152 = io_br_stall ? valid_99 : _GEN_1381; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2153 = io_br_stall ? valid_100 : _GEN_1382; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2154 = io_br_stall ? valid_101 : _GEN_1383; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2155 = io_br_stall ? valid_102 : _GEN_1384; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2156 = io_br_stall ? valid_103 : _GEN_1385; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2157 = io_br_stall ? valid_104 : _GEN_1386; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2158 = io_br_stall ? valid_105 : _GEN_1387; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2159 = io_br_stall ? valid_106 : _GEN_1388; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2160 = io_br_stall ? valid_107 : _GEN_1389; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2161 = io_br_stall ? valid_108 : _GEN_1390; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2162 = io_br_stall ? valid_109 : _GEN_1391; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2163 = io_br_stall ? valid_110 : _GEN_1392; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2164 = io_br_stall ? valid_111 : _GEN_1393; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2165 = io_br_stall ? valid_112 : _GEN_1394; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2166 = io_br_stall ? valid_113 : _GEN_1395; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2167 = io_br_stall ? valid_114 : _GEN_1396; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2168 = io_br_stall ? valid_115 : _GEN_1397; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2169 = io_br_stall ? valid_116 : _GEN_1398; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2170 = io_br_stall ? valid_117 : _GEN_1399; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2171 = io_br_stall ? valid_118 : _GEN_1400; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2172 = io_br_stall ? valid_119 : _GEN_1401; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2173 = io_br_stall ? valid_120 : _GEN_1402; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2174 = io_br_stall ? valid_121 : _GEN_1403; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2175 = io_br_stall ? valid_122 : _GEN_1404; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2176 = io_br_stall ? valid_123 : _GEN_1405; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2177 = io_br_stall ? valid_124 : _GEN_1406; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2178 = io_br_stall ? valid_125 : _GEN_1407; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2179 = io_br_stall ? valid_126 : _GEN_1408; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2180 = io_br_stall ? valid_127 : _GEN_1409; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2181 = io_br_stall ? valid_128 : _GEN_1410; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2182 = io_br_stall ? valid_129 : _GEN_1411; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2183 = io_br_stall ? valid_130 : _GEN_1412; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2184 = io_br_stall ? valid_131 : _GEN_1413; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2185 = io_br_stall ? valid_132 : _GEN_1414; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2186 = io_br_stall ? valid_133 : _GEN_1415; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2187 = io_br_stall ? valid_134 : _GEN_1416; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2188 = io_br_stall ? valid_135 : _GEN_1417; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2189 = io_br_stall ? valid_136 : _GEN_1418; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2190 = io_br_stall ? valid_137 : _GEN_1419; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2191 = io_br_stall ? valid_138 : _GEN_1420; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2192 = io_br_stall ? valid_139 : _GEN_1421; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2193 = io_br_stall ? valid_140 : _GEN_1422; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2194 = io_br_stall ? valid_141 : _GEN_1423; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2195 = io_br_stall ? valid_142 : _GEN_1424; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2196 = io_br_stall ? valid_143 : _GEN_1425; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2197 = io_br_stall ? valid_144 : _GEN_1426; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2198 = io_br_stall ? valid_145 : _GEN_1427; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2199 = io_br_stall ? valid_146 : _GEN_1428; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2200 = io_br_stall ? valid_147 : _GEN_1429; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2201 = io_br_stall ? valid_148 : _GEN_1430; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2202 = io_br_stall ? valid_149 : _GEN_1431; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2203 = io_br_stall ? valid_150 : _GEN_1432; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2204 = io_br_stall ? valid_151 : _GEN_1433; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2205 = io_br_stall ? valid_152 : _GEN_1434; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2206 = io_br_stall ? valid_153 : _GEN_1435; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2207 = io_br_stall ? valid_154 : _GEN_1436; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2208 = io_br_stall ? valid_155 : _GEN_1437; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2209 = io_br_stall ? valid_156 : _GEN_1438; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2210 = io_br_stall ? valid_157 : _GEN_1439; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2211 = io_br_stall ? valid_158 : _GEN_1440; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2212 = io_br_stall ? valid_159 : _GEN_1441; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2213 = io_br_stall ? valid_160 : _GEN_1442; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2214 = io_br_stall ? valid_161 : _GEN_1443; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2215 = io_br_stall ? valid_162 : _GEN_1444; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2216 = io_br_stall ? valid_163 : _GEN_1445; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2217 = io_br_stall ? valid_164 : _GEN_1446; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2218 = io_br_stall ? valid_165 : _GEN_1447; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2219 = io_br_stall ? valid_166 : _GEN_1448; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2220 = io_br_stall ? valid_167 : _GEN_1449; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2221 = io_br_stall ? valid_168 : _GEN_1450; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2222 = io_br_stall ? valid_169 : _GEN_1451; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2223 = io_br_stall ? valid_170 : _GEN_1452; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2224 = io_br_stall ? valid_171 : _GEN_1453; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2225 = io_br_stall ? valid_172 : _GEN_1454; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2226 = io_br_stall ? valid_173 : _GEN_1455; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2227 = io_br_stall ? valid_174 : _GEN_1456; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2228 = io_br_stall ? valid_175 : _GEN_1457; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2229 = io_br_stall ? valid_176 : _GEN_1458; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2230 = io_br_stall ? valid_177 : _GEN_1459; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2231 = io_br_stall ? valid_178 : _GEN_1460; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2232 = io_br_stall ? valid_179 : _GEN_1461; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2233 = io_br_stall ? valid_180 : _GEN_1462; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2234 = io_br_stall ? valid_181 : _GEN_1463; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2235 = io_br_stall ? valid_182 : _GEN_1464; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2236 = io_br_stall ? valid_183 : _GEN_1465; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2237 = io_br_stall ? valid_184 : _GEN_1466; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2238 = io_br_stall ? valid_185 : _GEN_1467; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2239 = io_br_stall ? valid_186 : _GEN_1468; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2240 = io_br_stall ? valid_187 : _GEN_1469; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2241 = io_br_stall ? valid_188 : _GEN_1470; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2242 = io_br_stall ? valid_189 : _GEN_1471; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2243 = io_br_stall ? valid_190 : _GEN_1472; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2244 = io_br_stall ? valid_191 : _GEN_1473; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2245 = io_br_stall ? valid_192 : _GEN_1474; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2246 = io_br_stall ? valid_193 : _GEN_1475; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2247 = io_br_stall ? valid_194 : _GEN_1476; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2248 = io_br_stall ? valid_195 : _GEN_1477; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2249 = io_br_stall ? valid_196 : _GEN_1478; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2250 = io_br_stall ? valid_197 : _GEN_1479; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2251 = io_br_stall ? valid_198 : _GEN_1480; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2252 = io_br_stall ? valid_199 : _GEN_1481; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2253 = io_br_stall ? valid_200 : _GEN_1482; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2254 = io_br_stall ? valid_201 : _GEN_1483; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2255 = io_br_stall ? valid_202 : _GEN_1484; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2256 = io_br_stall ? valid_203 : _GEN_1485; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2257 = io_br_stall ? valid_204 : _GEN_1486; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2258 = io_br_stall ? valid_205 : _GEN_1487; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2259 = io_br_stall ? valid_206 : _GEN_1488; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2260 = io_br_stall ? valid_207 : _GEN_1489; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2261 = io_br_stall ? valid_208 : _GEN_1490; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2262 = io_br_stall ? valid_209 : _GEN_1491; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2263 = io_br_stall ? valid_210 : _GEN_1492; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2264 = io_br_stall ? valid_211 : _GEN_1493; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2265 = io_br_stall ? valid_212 : _GEN_1494; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2266 = io_br_stall ? valid_213 : _GEN_1495; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2267 = io_br_stall ? valid_214 : _GEN_1496; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2268 = io_br_stall ? valid_215 : _GEN_1497; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2269 = io_br_stall ? valid_216 : _GEN_1498; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2270 = io_br_stall ? valid_217 : _GEN_1499; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2271 = io_br_stall ? valid_218 : _GEN_1500; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2272 = io_br_stall ? valid_219 : _GEN_1501; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2273 = io_br_stall ? valid_220 : _GEN_1502; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2274 = io_br_stall ? valid_221 : _GEN_1503; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2275 = io_br_stall ? valid_222 : _GEN_1504; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2276 = io_br_stall ? valid_223 : _GEN_1505; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2277 = io_br_stall ? valid_224 : _GEN_1506; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2278 = io_br_stall ? valid_225 : _GEN_1507; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2279 = io_br_stall ? valid_226 : _GEN_1508; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2280 = io_br_stall ? valid_227 : _GEN_1509; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2281 = io_br_stall ? valid_228 : _GEN_1510; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2282 = io_br_stall ? valid_229 : _GEN_1511; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2283 = io_br_stall ? valid_230 : _GEN_1512; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2284 = io_br_stall ? valid_231 : _GEN_1513; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2285 = io_br_stall ? valid_232 : _GEN_1514; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2286 = io_br_stall ? valid_233 : _GEN_1515; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2287 = io_br_stall ? valid_234 : _GEN_1516; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2288 = io_br_stall ? valid_235 : _GEN_1517; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2289 = io_br_stall ? valid_236 : _GEN_1518; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2290 = io_br_stall ? valid_237 : _GEN_1519; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2291 = io_br_stall ? valid_238 : _GEN_1520; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2292 = io_br_stall ? valid_239 : _GEN_1521; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2293 = io_br_stall ? valid_240 : _GEN_1522; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2294 = io_br_stall ? valid_241 : _GEN_1523; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2295 = io_br_stall ? valid_242 : _GEN_1524; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2296 = io_br_stall ? valid_243 : _GEN_1525; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2297 = io_br_stall ? valid_244 : _GEN_1526; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2298 = io_br_stall ? valid_245 : _GEN_1527; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2299 = io_br_stall ? valid_246 : _GEN_1528; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2300 = io_br_stall ? valid_247 : _GEN_1529; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2301 = io_br_stall ? valid_248 : _GEN_1530; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2302 = io_br_stall ? valid_249 : _GEN_1531; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2303 = io_br_stall ? valid_250 : _GEN_1532; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2304 = io_br_stall ? valid_251 : _GEN_1533; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2305 = io_br_stall ? valid_252 : _GEN_1534; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2306 = io_br_stall ? valid_253 : _GEN_1535; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2307 = io_br_stall ? valid_254 : _GEN_1536; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire  _GEN_2308 = io_br_stall ? valid_255 : _GEN_1537; // @[Icache.scala 73:26 Icache.scala 18:24]
  wire [19:0] _GEN_2309 = io_br_stall ? tag_0 : _GEN_1538; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2310 = io_br_stall ? tag_1 : _GEN_1539; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2311 = io_br_stall ? tag_2 : _GEN_1540; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2312 = io_br_stall ? tag_3 : _GEN_1541; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2313 = io_br_stall ? tag_4 : _GEN_1542; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2314 = io_br_stall ? tag_5 : _GEN_1543; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2315 = io_br_stall ? tag_6 : _GEN_1544; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2316 = io_br_stall ? tag_7 : _GEN_1545; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2317 = io_br_stall ? tag_8 : _GEN_1546; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2318 = io_br_stall ? tag_9 : _GEN_1547; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2319 = io_br_stall ? tag_10 : _GEN_1548; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2320 = io_br_stall ? tag_11 : _GEN_1549; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2321 = io_br_stall ? tag_12 : _GEN_1550; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2322 = io_br_stall ? tag_13 : _GEN_1551; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2323 = io_br_stall ? tag_14 : _GEN_1552; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2324 = io_br_stall ? tag_15 : _GEN_1553; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2325 = io_br_stall ? tag_16 : _GEN_1554; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2326 = io_br_stall ? tag_17 : _GEN_1555; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2327 = io_br_stall ? tag_18 : _GEN_1556; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2328 = io_br_stall ? tag_19 : _GEN_1557; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2329 = io_br_stall ? tag_20 : _GEN_1558; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2330 = io_br_stall ? tag_21 : _GEN_1559; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2331 = io_br_stall ? tag_22 : _GEN_1560; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2332 = io_br_stall ? tag_23 : _GEN_1561; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2333 = io_br_stall ? tag_24 : _GEN_1562; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2334 = io_br_stall ? tag_25 : _GEN_1563; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2335 = io_br_stall ? tag_26 : _GEN_1564; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2336 = io_br_stall ? tag_27 : _GEN_1565; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2337 = io_br_stall ? tag_28 : _GEN_1566; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2338 = io_br_stall ? tag_29 : _GEN_1567; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2339 = io_br_stall ? tag_30 : _GEN_1568; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2340 = io_br_stall ? tag_31 : _GEN_1569; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2341 = io_br_stall ? tag_32 : _GEN_1570; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2342 = io_br_stall ? tag_33 : _GEN_1571; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2343 = io_br_stall ? tag_34 : _GEN_1572; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2344 = io_br_stall ? tag_35 : _GEN_1573; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2345 = io_br_stall ? tag_36 : _GEN_1574; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2346 = io_br_stall ? tag_37 : _GEN_1575; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2347 = io_br_stall ? tag_38 : _GEN_1576; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2348 = io_br_stall ? tag_39 : _GEN_1577; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2349 = io_br_stall ? tag_40 : _GEN_1578; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2350 = io_br_stall ? tag_41 : _GEN_1579; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2351 = io_br_stall ? tag_42 : _GEN_1580; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2352 = io_br_stall ? tag_43 : _GEN_1581; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2353 = io_br_stall ? tag_44 : _GEN_1582; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2354 = io_br_stall ? tag_45 : _GEN_1583; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2355 = io_br_stall ? tag_46 : _GEN_1584; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2356 = io_br_stall ? tag_47 : _GEN_1585; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2357 = io_br_stall ? tag_48 : _GEN_1586; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2358 = io_br_stall ? tag_49 : _GEN_1587; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2359 = io_br_stall ? tag_50 : _GEN_1588; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2360 = io_br_stall ? tag_51 : _GEN_1589; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2361 = io_br_stall ? tag_52 : _GEN_1590; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2362 = io_br_stall ? tag_53 : _GEN_1591; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2363 = io_br_stall ? tag_54 : _GEN_1592; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2364 = io_br_stall ? tag_55 : _GEN_1593; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2365 = io_br_stall ? tag_56 : _GEN_1594; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2366 = io_br_stall ? tag_57 : _GEN_1595; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2367 = io_br_stall ? tag_58 : _GEN_1596; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2368 = io_br_stall ? tag_59 : _GEN_1597; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2369 = io_br_stall ? tag_60 : _GEN_1598; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2370 = io_br_stall ? tag_61 : _GEN_1599; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2371 = io_br_stall ? tag_62 : _GEN_1600; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2372 = io_br_stall ? tag_63 : _GEN_1601; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2373 = io_br_stall ? tag_64 : _GEN_1602; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2374 = io_br_stall ? tag_65 : _GEN_1603; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2375 = io_br_stall ? tag_66 : _GEN_1604; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2376 = io_br_stall ? tag_67 : _GEN_1605; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2377 = io_br_stall ? tag_68 : _GEN_1606; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2378 = io_br_stall ? tag_69 : _GEN_1607; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2379 = io_br_stall ? tag_70 : _GEN_1608; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2380 = io_br_stall ? tag_71 : _GEN_1609; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2381 = io_br_stall ? tag_72 : _GEN_1610; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2382 = io_br_stall ? tag_73 : _GEN_1611; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2383 = io_br_stall ? tag_74 : _GEN_1612; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2384 = io_br_stall ? tag_75 : _GEN_1613; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2385 = io_br_stall ? tag_76 : _GEN_1614; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2386 = io_br_stall ? tag_77 : _GEN_1615; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2387 = io_br_stall ? tag_78 : _GEN_1616; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2388 = io_br_stall ? tag_79 : _GEN_1617; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2389 = io_br_stall ? tag_80 : _GEN_1618; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2390 = io_br_stall ? tag_81 : _GEN_1619; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2391 = io_br_stall ? tag_82 : _GEN_1620; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2392 = io_br_stall ? tag_83 : _GEN_1621; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2393 = io_br_stall ? tag_84 : _GEN_1622; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2394 = io_br_stall ? tag_85 : _GEN_1623; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2395 = io_br_stall ? tag_86 : _GEN_1624; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2396 = io_br_stall ? tag_87 : _GEN_1625; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2397 = io_br_stall ? tag_88 : _GEN_1626; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2398 = io_br_stall ? tag_89 : _GEN_1627; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2399 = io_br_stall ? tag_90 : _GEN_1628; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2400 = io_br_stall ? tag_91 : _GEN_1629; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2401 = io_br_stall ? tag_92 : _GEN_1630; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2402 = io_br_stall ? tag_93 : _GEN_1631; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2403 = io_br_stall ? tag_94 : _GEN_1632; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2404 = io_br_stall ? tag_95 : _GEN_1633; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2405 = io_br_stall ? tag_96 : _GEN_1634; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2406 = io_br_stall ? tag_97 : _GEN_1635; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2407 = io_br_stall ? tag_98 : _GEN_1636; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2408 = io_br_stall ? tag_99 : _GEN_1637; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2409 = io_br_stall ? tag_100 : _GEN_1638; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2410 = io_br_stall ? tag_101 : _GEN_1639; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2411 = io_br_stall ? tag_102 : _GEN_1640; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2412 = io_br_stall ? tag_103 : _GEN_1641; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2413 = io_br_stall ? tag_104 : _GEN_1642; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2414 = io_br_stall ? tag_105 : _GEN_1643; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2415 = io_br_stall ? tag_106 : _GEN_1644; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2416 = io_br_stall ? tag_107 : _GEN_1645; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2417 = io_br_stall ? tag_108 : _GEN_1646; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2418 = io_br_stall ? tag_109 : _GEN_1647; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2419 = io_br_stall ? tag_110 : _GEN_1648; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2420 = io_br_stall ? tag_111 : _GEN_1649; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2421 = io_br_stall ? tag_112 : _GEN_1650; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2422 = io_br_stall ? tag_113 : _GEN_1651; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2423 = io_br_stall ? tag_114 : _GEN_1652; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2424 = io_br_stall ? tag_115 : _GEN_1653; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2425 = io_br_stall ? tag_116 : _GEN_1654; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2426 = io_br_stall ? tag_117 : _GEN_1655; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2427 = io_br_stall ? tag_118 : _GEN_1656; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2428 = io_br_stall ? tag_119 : _GEN_1657; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2429 = io_br_stall ? tag_120 : _GEN_1658; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2430 = io_br_stall ? tag_121 : _GEN_1659; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2431 = io_br_stall ? tag_122 : _GEN_1660; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2432 = io_br_stall ? tag_123 : _GEN_1661; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2433 = io_br_stall ? tag_124 : _GEN_1662; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2434 = io_br_stall ? tag_125 : _GEN_1663; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2435 = io_br_stall ? tag_126 : _GEN_1664; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2436 = io_br_stall ? tag_127 : _GEN_1665; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2437 = io_br_stall ? tag_128 : _GEN_1666; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2438 = io_br_stall ? tag_129 : _GEN_1667; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2439 = io_br_stall ? tag_130 : _GEN_1668; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2440 = io_br_stall ? tag_131 : _GEN_1669; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2441 = io_br_stall ? tag_132 : _GEN_1670; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2442 = io_br_stall ? tag_133 : _GEN_1671; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2443 = io_br_stall ? tag_134 : _GEN_1672; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2444 = io_br_stall ? tag_135 : _GEN_1673; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2445 = io_br_stall ? tag_136 : _GEN_1674; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2446 = io_br_stall ? tag_137 : _GEN_1675; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2447 = io_br_stall ? tag_138 : _GEN_1676; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2448 = io_br_stall ? tag_139 : _GEN_1677; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2449 = io_br_stall ? tag_140 : _GEN_1678; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2450 = io_br_stall ? tag_141 : _GEN_1679; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2451 = io_br_stall ? tag_142 : _GEN_1680; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2452 = io_br_stall ? tag_143 : _GEN_1681; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2453 = io_br_stall ? tag_144 : _GEN_1682; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2454 = io_br_stall ? tag_145 : _GEN_1683; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2455 = io_br_stall ? tag_146 : _GEN_1684; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2456 = io_br_stall ? tag_147 : _GEN_1685; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2457 = io_br_stall ? tag_148 : _GEN_1686; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2458 = io_br_stall ? tag_149 : _GEN_1687; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2459 = io_br_stall ? tag_150 : _GEN_1688; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2460 = io_br_stall ? tag_151 : _GEN_1689; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2461 = io_br_stall ? tag_152 : _GEN_1690; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2462 = io_br_stall ? tag_153 : _GEN_1691; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2463 = io_br_stall ? tag_154 : _GEN_1692; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2464 = io_br_stall ? tag_155 : _GEN_1693; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2465 = io_br_stall ? tag_156 : _GEN_1694; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2466 = io_br_stall ? tag_157 : _GEN_1695; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2467 = io_br_stall ? tag_158 : _GEN_1696; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2468 = io_br_stall ? tag_159 : _GEN_1697; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2469 = io_br_stall ? tag_160 : _GEN_1698; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2470 = io_br_stall ? tag_161 : _GEN_1699; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2471 = io_br_stall ? tag_162 : _GEN_1700; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2472 = io_br_stall ? tag_163 : _GEN_1701; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2473 = io_br_stall ? tag_164 : _GEN_1702; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2474 = io_br_stall ? tag_165 : _GEN_1703; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2475 = io_br_stall ? tag_166 : _GEN_1704; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2476 = io_br_stall ? tag_167 : _GEN_1705; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2477 = io_br_stall ? tag_168 : _GEN_1706; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2478 = io_br_stall ? tag_169 : _GEN_1707; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2479 = io_br_stall ? tag_170 : _GEN_1708; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2480 = io_br_stall ? tag_171 : _GEN_1709; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2481 = io_br_stall ? tag_172 : _GEN_1710; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2482 = io_br_stall ? tag_173 : _GEN_1711; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2483 = io_br_stall ? tag_174 : _GEN_1712; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2484 = io_br_stall ? tag_175 : _GEN_1713; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2485 = io_br_stall ? tag_176 : _GEN_1714; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2486 = io_br_stall ? tag_177 : _GEN_1715; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2487 = io_br_stall ? tag_178 : _GEN_1716; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2488 = io_br_stall ? tag_179 : _GEN_1717; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2489 = io_br_stall ? tag_180 : _GEN_1718; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2490 = io_br_stall ? tag_181 : _GEN_1719; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2491 = io_br_stall ? tag_182 : _GEN_1720; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2492 = io_br_stall ? tag_183 : _GEN_1721; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2493 = io_br_stall ? tag_184 : _GEN_1722; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2494 = io_br_stall ? tag_185 : _GEN_1723; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2495 = io_br_stall ? tag_186 : _GEN_1724; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2496 = io_br_stall ? tag_187 : _GEN_1725; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2497 = io_br_stall ? tag_188 : _GEN_1726; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2498 = io_br_stall ? tag_189 : _GEN_1727; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2499 = io_br_stall ? tag_190 : _GEN_1728; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2500 = io_br_stall ? tag_191 : _GEN_1729; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2501 = io_br_stall ? tag_192 : _GEN_1730; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2502 = io_br_stall ? tag_193 : _GEN_1731; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2503 = io_br_stall ? tag_194 : _GEN_1732; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2504 = io_br_stall ? tag_195 : _GEN_1733; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2505 = io_br_stall ? tag_196 : _GEN_1734; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2506 = io_br_stall ? tag_197 : _GEN_1735; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2507 = io_br_stall ? tag_198 : _GEN_1736; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2508 = io_br_stall ? tag_199 : _GEN_1737; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2509 = io_br_stall ? tag_200 : _GEN_1738; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2510 = io_br_stall ? tag_201 : _GEN_1739; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2511 = io_br_stall ? tag_202 : _GEN_1740; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2512 = io_br_stall ? tag_203 : _GEN_1741; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2513 = io_br_stall ? tag_204 : _GEN_1742; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2514 = io_br_stall ? tag_205 : _GEN_1743; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2515 = io_br_stall ? tag_206 : _GEN_1744; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2516 = io_br_stall ? tag_207 : _GEN_1745; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2517 = io_br_stall ? tag_208 : _GEN_1746; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2518 = io_br_stall ? tag_209 : _GEN_1747; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2519 = io_br_stall ? tag_210 : _GEN_1748; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2520 = io_br_stall ? tag_211 : _GEN_1749; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2521 = io_br_stall ? tag_212 : _GEN_1750; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2522 = io_br_stall ? tag_213 : _GEN_1751; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2523 = io_br_stall ? tag_214 : _GEN_1752; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2524 = io_br_stall ? tag_215 : _GEN_1753; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2525 = io_br_stall ? tag_216 : _GEN_1754; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2526 = io_br_stall ? tag_217 : _GEN_1755; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2527 = io_br_stall ? tag_218 : _GEN_1756; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2528 = io_br_stall ? tag_219 : _GEN_1757; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2529 = io_br_stall ? tag_220 : _GEN_1758; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2530 = io_br_stall ? tag_221 : _GEN_1759; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2531 = io_br_stall ? tag_222 : _GEN_1760; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2532 = io_br_stall ? tag_223 : _GEN_1761; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2533 = io_br_stall ? tag_224 : _GEN_1762; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2534 = io_br_stall ? tag_225 : _GEN_1763; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2535 = io_br_stall ? tag_226 : _GEN_1764; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2536 = io_br_stall ? tag_227 : _GEN_1765; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2537 = io_br_stall ? tag_228 : _GEN_1766; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2538 = io_br_stall ? tag_229 : _GEN_1767; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2539 = io_br_stall ? tag_230 : _GEN_1768; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2540 = io_br_stall ? tag_231 : _GEN_1769; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2541 = io_br_stall ? tag_232 : _GEN_1770; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2542 = io_br_stall ? tag_233 : _GEN_1771; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2543 = io_br_stall ? tag_234 : _GEN_1772; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2544 = io_br_stall ? tag_235 : _GEN_1773; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2545 = io_br_stall ? tag_236 : _GEN_1774; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2546 = io_br_stall ? tag_237 : _GEN_1775; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2547 = io_br_stall ? tag_238 : _GEN_1776; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2548 = io_br_stall ? tag_239 : _GEN_1777; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2549 = io_br_stall ? tag_240 : _GEN_1778; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2550 = io_br_stall ? tag_241 : _GEN_1779; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2551 = io_br_stall ? tag_242 : _GEN_1780; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2552 = io_br_stall ? tag_243 : _GEN_1781; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2553 = io_br_stall ? tag_244 : _GEN_1782; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2554 = io_br_stall ? tag_245 : _GEN_1783; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2555 = io_br_stall ? tag_246 : _GEN_1784; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2556 = io_br_stall ? tag_247 : _GEN_1785; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2557 = io_br_stall ? tag_248 : _GEN_1786; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2558 = io_br_stall ? tag_249 : _GEN_1787; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2559 = io_br_stall ? tag_250 : _GEN_1788; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2560 = io_br_stall ? tag_251 : _GEN_1789; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2561 = io_br_stall ? tag_252 : _GEN_1790; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2562 = io_br_stall ? tag_253 : _GEN_1791; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2563 = io_br_stall ? tag_254 : _GEN_1792; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire [19:0] _GEN_2564 = io_br_stall ? tag_255 : _GEN_1793; // @[Icache.scala 73:26 Icache.scala 17:24]
  wire  _GEN_2821 = io_br_stall ? inst_ready : _GEN_2050; // @[Icache.scala 73:26 Icache.scala 42:28]
  wire  _T_3 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = ~cache_fill; // @[Icache.scala 89:13]
  wire [2:0] _GEN_2822 = ~cache_fill ? 3'h3 : 3'h4; // @[Icache.scala 89:26 Icache.scala 90:15 Icache.scala 97:15]
  wire [31:0] _GEN_2825 = ~cache_fill ? io_imem_inst_addr : 32'h0; // @[Icache.scala 89:26 Icache.scala 93:21]
  wire  _GEN_2827 = io_out_inst_ready | cache_fill; // @[Icache.scala 99:29 Icache.scala 100:21 Icache.scala 51:28]
  wire  _GEN_2828 = io_out_inst_ready | cache_wen; // @[Icache.scala 99:29 Icache.scala 101:21 Icache.scala 52:28]
  wire [127:0] _GEN_2829 = io_out_inst_ready ? io_out_inst_read : cache_wdata; // @[Icache.scala 99:29 Icache.scala 102:21 Icache.scala 53:28]
  wire  _GEN_2830 = io_out_inst_ready ? 1'h0 : _T_4; // @[Icache.scala 99:29 Icache.scala 103:21]
  wire  _T_5 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _GEN_3599 = _T_5 ? 1'h0 : cache_fill; // @[Conditional.scala 39:67 Icache.scala 108:25 Icache.scala 51:28]
  wire  _GEN_3600 = _T_5 | inst_ready; // @[Conditional.scala 39:67 Icache.scala 109:25 Icache.scala 42:28]
  wire  _GEN_3601 = _T_5 ? 1'h0 : cache_wen; // @[Conditional.scala 39:67 Icache.scala 110:25 Icache.scala 52:28]
  wire  _GEN_3602 = _T_5 ? _GEN_514 : valid_0; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3603 = _T_5 ? _GEN_515 : valid_1; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3604 = _T_5 ? _GEN_516 : valid_2; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3605 = _T_5 ? _GEN_517 : valid_3; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3606 = _T_5 ? _GEN_518 : valid_4; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3607 = _T_5 ? _GEN_519 : valid_5; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3608 = _T_5 ? _GEN_520 : valid_6; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3609 = _T_5 ? _GEN_521 : valid_7; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3610 = _T_5 ? _GEN_522 : valid_8; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3611 = _T_5 ? _GEN_523 : valid_9; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3612 = _T_5 ? _GEN_524 : valid_10; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3613 = _T_5 ? _GEN_525 : valid_11; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3614 = _T_5 ? _GEN_526 : valid_12; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3615 = _T_5 ? _GEN_527 : valid_13; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3616 = _T_5 ? _GEN_528 : valid_14; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3617 = _T_5 ? _GEN_529 : valid_15; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3618 = _T_5 ? _GEN_530 : valid_16; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3619 = _T_5 ? _GEN_531 : valid_17; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3620 = _T_5 ? _GEN_532 : valid_18; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3621 = _T_5 ? _GEN_533 : valid_19; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3622 = _T_5 ? _GEN_534 : valid_20; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3623 = _T_5 ? _GEN_535 : valid_21; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3624 = _T_5 ? _GEN_536 : valid_22; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3625 = _T_5 ? _GEN_537 : valid_23; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3626 = _T_5 ? _GEN_538 : valid_24; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3627 = _T_5 ? _GEN_539 : valid_25; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3628 = _T_5 ? _GEN_540 : valid_26; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3629 = _T_5 ? _GEN_541 : valid_27; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3630 = _T_5 ? _GEN_542 : valid_28; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3631 = _T_5 ? _GEN_543 : valid_29; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3632 = _T_5 ? _GEN_544 : valid_30; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3633 = _T_5 ? _GEN_545 : valid_31; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3634 = _T_5 ? _GEN_546 : valid_32; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3635 = _T_5 ? _GEN_547 : valid_33; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3636 = _T_5 ? _GEN_548 : valid_34; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3637 = _T_5 ? _GEN_549 : valid_35; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3638 = _T_5 ? _GEN_550 : valid_36; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3639 = _T_5 ? _GEN_551 : valid_37; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3640 = _T_5 ? _GEN_552 : valid_38; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3641 = _T_5 ? _GEN_553 : valid_39; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3642 = _T_5 ? _GEN_554 : valid_40; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3643 = _T_5 ? _GEN_555 : valid_41; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3644 = _T_5 ? _GEN_556 : valid_42; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3645 = _T_5 ? _GEN_557 : valid_43; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3646 = _T_5 ? _GEN_558 : valid_44; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3647 = _T_5 ? _GEN_559 : valid_45; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3648 = _T_5 ? _GEN_560 : valid_46; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3649 = _T_5 ? _GEN_561 : valid_47; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3650 = _T_5 ? _GEN_562 : valid_48; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3651 = _T_5 ? _GEN_563 : valid_49; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3652 = _T_5 ? _GEN_564 : valid_50; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3653 = _T_5 ? _GEN_565 : valid_51; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3654 = _T_5 ? _GEN_566 : valid_52; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3655 = _T_5 ? _GEN_567 : valid_53; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3656 = _T_5 ? _GEN_568 : valid_54; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3657 = _T_5 ? _GEN_569 : valid_55; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3658 = _T_5 ? _GEN_570 : valid_56; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3659 = _T_5 ? _GEN_571 : valid_57; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3660 = _T_5 ? _GEN_572 : valid_58; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3661 = _T_5 ? _GEN_573 : valid_59; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3662 = _T_5 ? _GEN_574 : valid_60; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3663 = _T_5 ? _GEN_575 : valid_61; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3664 = _T_5 ? _GEN_576 : valid_62; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3665 = _T_5 ? _GEN_577 : valid_63; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3666 = _T_5 ? _GEN_578 : valid_64; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3667 = _T_5 ? _GEN_579 : valid_65; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3668 = _T_5 ? _GEN_580 : valid_66; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3669 = _T_5 ? _GEN_581 : valid_67; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3670 = _T_5 ? _GEN_582 : valid_68; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3671 = _T_5 ? _GEN_583 : valid_69; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3672 = _T_5 ? _GEN_584 : valid_70; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3673 = _T_5 ? _GEN_585 : valid_71; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3674 = _T_5 ? _GEN_586 : valid_72; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3675 = _T_5 ? _GEN_587 : valid_73; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3676 = _T_5 ? _GEN_588 : valid_74; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3677 = _T_5 ? _GEN_589 : valid_75; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3678 = _T_5 ? _GEN_590 : valid_76; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3679 = _T_5 ? _GEN_591 : valid_77; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3680 = _T_5 ? _GEN_592 : valid_78; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3681 = _T_5 ? _GEN_593 : valid_79; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3682 = _T_5 ? _GEN_594 : valid_80; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3683 = _T_5 ? _GEN_595 : valid_81; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3684 = _T_5 ? _GEN_596 : valid_82; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3685 = _T_5 ? _GEN_597 : valid_83; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3686 = _T_5 ? _GEN_598 : valid_84; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3687 = _T_5 ? _GEN_599 : valid_85; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3688 = _T_5 ? _GEN_600 : valid_86; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3689 = _T_5 ? _GEN_601 : valid_87; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3690 = _T_5 ? _GEN_602 : valid_88; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3691 = _T_5 ? _GEN_603 : valid_89; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3692 = _T_5 ? _GEN_604 : valid_90; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3693 = _T_5 ? _GEN_605 : valid_91; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3694 = _T_5 ? _GEN_606 : valid_92; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3695 = _T_5 ? _GEN_607 : valid_93; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3696 = _T_5 ? _GEN_608 : valid_94; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3697 = _T_5 ? _GEN_609 : valid_95; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3698 = _T_5 ? _GEN_610 : valid_96; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3699 = _T_5 ? _GEN_611 : valid_97; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3700 = _T_5 ? _GEN_612 : valid_98; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3701 = _T_5 ? _GEN_613 : valid_99; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3702 = _T_5 ? _GEN_614 : valid_100; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3703 = _T_5 ? _GEN_615 : valid_101; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3704 = _T_5 ? _GEN_616 : valid_102; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3705 = _T_5 ? _GEN_617 : valid_103; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3706 = _T_5 ? _GEN_618 : valid_104; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3707 = _T_5 ? _GEN_619 : valid_105; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3708 = _T_5 ? _GEN_620 : valid_106; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3709 = _T_5 ? _GEN_621 : valid_107; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3710 = _T_5 ? _GEN_622 : valid_108; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3711 = _T_5 ? _GEN_623 : valid_109; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3712 = _T_5 ? _GEN_624 : valid_110; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3713 = _T_5 ? _GEN_625 : valid_111; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3714 = _T_5 ? _GEN_626 : valid_112; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3715 = _T_5 ? _GEN_627 : valid_113; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3716 = _T_5 ? _GEN_628 : valid_114; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3717 = _T_5 ? _GEN_629 : valid_115; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3718 = _T_5 ? _GEN_630 : valid_116; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3719 = _T_5 ? _GEN_631 : valid_117; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3720 = _T_5 ? _GEN_632 : valid_118; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3721 = _T_5 ? _GEN_633 : valid_119; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3722 = _T_5 ? _GEN_634 : valid_120; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3723 = _T_5 ? _GEN_635 : valid_121; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3724 = _T_5 ? _GEN_636 : valid_122; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3725 = _T_5 ? _GEN_637 : valid_123; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3726 = _T_5 ? _GEN_638 : valid_124; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3727 = _T_5 ? _GEN_639 : valid_125; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3728 = _T_5 ? _GEN_640 : valid_126; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3729 = _T_5 ? _GEN_641 : valid_127; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3730 = _T_5 ? _GEN_642 : valid_128; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3731 = _T_5 ? _GEN_643 : valid_129; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3732 = _T_5 ? _GEN_644 : valid_130; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3733 = _T_5 ? _GEN_645 : valid_131; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3734 = _T_5 ? _GEN_646 : valid_132; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3735 = _T_5 ? _GEN_647 : valid_133; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3736 = _T_5 ? _GEN_648 : valid_134; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3737 = _T_5 ? _GEN_649 : valid_135; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3738 = _T_5 ? _GEN_650 : valid_136; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3739 = _T_5 ? _GEN_651 : valid_137; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3740 = _T_5 ? _GEN_652 : valid_138; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3741 = _T_5 ? _GEN_653 : valid_139; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3742 = _T_5 ? _GEN_654 : valid_140; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3743 = _T_5 ? _GEN_655 : valid_141; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3744 = _T_5 ? _GEN_656 : valid_142; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3745 = _T_5 ? _GEN_657 : valid_143; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3746 = _T_5 ? _GEN_658 : valid_144; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3747 = _T_5 ? _GEN_659 : valid_145; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3748 = _T_5 ? _GEN_660 : valid_146; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3749 = _T_5 ? _GEN_661 : valid_147; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3750 = _T_5 ? _GEN_662 : valid_148; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3751 = _T_5 ? _GEN_663 : valid_149; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3752 = _T_5 ? _GEN_664 : valid_150; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3753 = _T_5 ? _GEN_665 : valid_151; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3754 = _T_5 ? _GEN_666 : valid_152; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3755 = _T_5 ? _GEN_667 : valid_153; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3756 = _T_5 ? _GEN_668 : valid_154; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3757 = _T_5 ? _GEN_669 : valid_155; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3758 = _T_5 ? _GEN_670 : valid_156; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3759 = _T_5 ? _GEN_671 : valid_157; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3760 = _T_5 ? _GEN_672 : valid_158; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3761 = _T_5 ? _GEN_673 : valid_159; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3762 = _T_5 ? _GEN_674 : valid_160; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3763 = _T_5 ? _GEN_675 : valid_161; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3764 = _T_5 ? _GEN_676 : valid_162; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3765 = _T_5 ? _GEN_677 : valid_163; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3766 = _T_5 ? _GEN_678 : valid_164; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3767 = _T_5 ? _GEN_679 : valid_165; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3768 = _T_5 ? _GEN_680 : valid_166; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3769 = _T_5 ? _GEN_681 : valid_167; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3770 = _T_5 ? _GEN_682 : valid_168; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3771 = _T_5 ? _GEN_683 : valid_169; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3772 = _T_5 ? _GEN_684 : valid_170; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3773 = _T_5 ? _GEN_685 : valid_171; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3774 = _T_5 ? _GEN_686 : valid_172; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3775 = _T_5 ? _GEN_687 : valid_173; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3776 = _T_5 ? _GEN_688 : valid_174; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3777 = _T_5 ? _GEN_689 : valid_175; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3778 = _T_5 ? _GEN_690 : valid_176; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3779 = _T_5 ? _GEN_691 : valid_177; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3780 = _T_5 ? _GEN_692 : valid_178; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3781 = _T_5 ? _GEN_693 : valid_179; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3782 = _T_5 ? _GEN_694 : valid_180; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3783 = _T_5 ? _GEN_695 : valid_181; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3784 = _T_5 ? _GEN_696 : valid_182; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3785 = _T_5 ? _GEN_697 : valid_183; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3786 = _T_5 ? _GEN_698 : valid_184; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3787 = _T_5 ? _GEN_699 : valid_185; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3788 = _T_5 ? _GEN_700 : valid_186; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3789 = _T_5 ? _GEN_701 : valid_187; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3790 = _T_5 ? _GEN_702 : valid_188; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3791 = _T_5 ? _GEN_703 : valid_189; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3792 = _T_5 ? _GEN_704 : valid_190; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3793 = _T_5 ? _GEN_705 : valid_191; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3794 = _T_5 ? _GEN_706 : valid_192; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3795 = _T_5 ? _GEN_707 : valid_193; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3796 = _T_5 ? _GEN_708 : valid_194; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3797 = _T_5 ? _GEN_709 : valid_195; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3798 = _T_5 ? _GEN_710 : valid_196; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3799 = _T_5 ? _GEN_711 : valid_197; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3800 = _T_5 ? _GEN_712 : valid_198; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3801 = _T_5 ? _GEN_713 : valid_199; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3802 = _T_5 ? _GEN_714 : valid_200; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3803 = _T_5 ? _GEN_715 : valid_201; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3804 = _T_5 ? _GEN_716 : valid_202; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3805 = _T_5 ? _GEN_717 : valid_203; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3806 = _T_5 ? _GEN_718 : valid_204; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3807 = _T_5 ? _GEN_719 : valid_205; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3808 = _T_5 ? _GEN_720 : valid_206; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3809 = _T_5 ? _GEN_721 : valid_207; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3810 = _T_5 ? _GEN_722 : valid_208; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3811 = _T_5 ? _GEN_723 : valid_209; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3812 = _T_5 ? _GEN_724 : valid_210; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3813 = _T_5 ? _GEN_725 : valid_211; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3814 = _T_5 ? _GEN_726 : valid_212; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3815 = _T_5 ? _GEN_727 : valid_213; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3816 = _T_5 ? _GEN_728 : valid_214; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3817 = _T_5 ? _GEN_729 : valid_215; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3818 = _T_5 ? _GEN_730 : valid_216; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3819 = _T_5 ? _GEN_731 : valid_217; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3820 = _T_5 ? _GEN_732 : valid_218; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3821 = _T_5 ? _GEN_733 : valid_219; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3822 = _T_5 ? _GEN_734 : valid_220; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3823 = _T_5 ? _GEN_735 : valid_221; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3824 = _T_5 ? _GEN_736 : valid_222; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3825 = _T_5 ? _GEN_737 : valid_223; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3826 = _T_5 ? _GEN_738 : valid_224; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3827 = _T_5 ? _GEN_739 : valid_225; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3828 = _T_5 ? _GEN_740 : valid_226; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3829 = _T_5 ? _GEN_741 : valid_227; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3830 = _T_5 ? _GEN_742 : valid_228; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3831 = _T_5 ? _GEN_743 : valid_229; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3832 = _T_5 ? _GEN_744 : valid_230; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3833 = _T_5 ? _GEN_745 : valid_231; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3834 = _T_5 ? _GEN_746 : valid_232; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3835 = _T_5 ? _GEN_747 : valid_233; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3836 = _T_5 ? _GEN_748 : valid_234; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3837 = _T_5 ? _GEN_749 : valid_235; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3838 = _T_5 ? _GEN_750 : valid_236; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3839 = _T_5 ? _GEN_751 : valid_237; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3840 = _T_5 ? _GEN_752 : valid_238; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3841 = _T_5 ? _GEN_753 : valid_239; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3842 = _T_5 ? _GEN_754 : valid_240; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3843 = _T_5 ? _GEN_755 : valid_241; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3844 = _T_5 ? _GEN_756 : valid_242; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3845 = _T_5 ? _GEN_757 : valid_243; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3846 = _T_5 ? _GEN_758 : valid_244; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3847 = _T_5 ? _GEN_759 : valid_245; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3848 = _T_5 ? _GEN_760 : valid_246; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3849 = _T_5 ? _GEN_761 : valid_247; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3850 = _T_5 ? _GEN_762 : valid_248; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3851 = _T_5 ? _GEN_763 : valid_249; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3852 = _T_5 ? _GEN_764 : valid_250; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3853 = _T_5 ? _GEN_765 : valid_251; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3854 = _T_5 ? _GEN_766 : valid_252; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3855 = _T_5 ? _GEN_767 : valid_253; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3856 = _T_5 ? _GEN_768 : valid_254; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_3857 = _T_5 ? _GEN_769 : valid_255; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire [19:0] _GEN_3858 = _T_5 ? _GEN_770 : tag_0; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3859 = _T_5 ? _GEN_771 : tag_1; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3860 = _T_5 ? _GEN_772 : tag_2; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3861 = _T_5 ? _GEN_773 : tag_3; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3862 = _T_5 ? _GEN_774 : tag_4; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3863 = _T_5 ? _GEN_775 : tag_5; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3864 = _T_5 ? _GEN_776 : tag_6; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3865 = _T_5 ? _GEN_777 : tag_7; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3866 = _T_5 ? _GEN_778 : tag_8; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3867 = _T_5 ? _GEN_779 : tag_9; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3868 = _T_5 ? _GEN_780 : tag_10; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3869 = _T_5 ? _GEN_781 : tag_11; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3870 = _T_5 ? _GEN_782 : tag_12; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3871 = _T_5 ? _GEN_783 : tag_13; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3872 = _T_5 ? _GEN_784 : tag_14; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3873 = _T_5 ? _GEN_785 : tag_15; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3874 = _T_5 ? _GEN_786 : tag_16; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3875 = _T_5 ? _GEN_787 : tag_17; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3876 = _T_5 ? _GEN_788 : tag_18; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3877 = _T_5 ? _GEN_789 : tag_19; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3878 = _T_5 ? _GEN_790 : tag_20; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3879 = _T_5 ? _GEN_791 : tag_21; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3880 = _T_5 ? _GEN_792 : tag_22; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3881 = _T_5 ? _GEN_793 : tag_23; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3882 = _T_5 ? _GEN_794 : tag_24; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3883 = _T_5 ? _GEN_795 : tag_25; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3884 = _T_5 ? _GEN_796 : tag_26; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3885 = _T_5 ? _GEN_797 : tag_27; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3886 = _T_5 ? _GEN_798 : tag_28; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3887 = _T_5 ? _GEN_799 : tag_29; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3888 = _T_5 ? _GEN_800 : tag_30; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3889 = _T_5 ? _GEN_801 : tag_31; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3890 = _T_5 ? _GEN_802 : tag_32; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3891 = _T_5 ? _GEN_803 : tag_33; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3892 = _T_5 ? _GEN_804 : tag_34; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3893 = _T_5 ? _GEN_805 : tag_35; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3894 = _T_5 ? _GEN_806 : tag_36; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3895 = _T_5 ? _GEN_807 : tag_37; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3896 = _T_5 ? _GEN_808 : tag_38; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3897 = _T_5 ? _GEN_809 : tag_39; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3898 = _T_5 ? _GEN_810 : tag_40; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3899 = _T_5 ? _GEN_811 : tag_41; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3900 = _T_5 ? _GEN_812 : tag_42; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3901 = _T_5 ? _GEN_813 : tag_43; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3902 = _T_5 ? _GEN_814 : tag_44; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3903 = _T_5 ? _GEN_815 : tag_45; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3904 = _T_5 ? _GEN_816 : tag_46; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3905 = _T_5 ? _GEN_817 : tag_47; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3906 = _T_5 ? _GEN_818 : tag_48; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3907 = _T_5 ? _GEN_819 : tag_49; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3908 = _T_5 ? _GEN_820 : tag_50; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3909 = _T_5 ? _GEN_821 : tag_51; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3910 = _T_5 ? _GEN_822 : tag_52; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3911 = _T_5 ? _GEN_823 : tag_53; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3912 = _T_5 ? _GEN_824 : tag_54; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3913 = _T_5 ? _GEN_825 : tag_55; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3914 = _T_5 ? _GEN_826 : tag_56; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3915 = _T_5 ? _GEN_827 : tag_57; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3916 = _T_5 ? _GEN_828 : tag_58; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3917 = _T_5 ? _GEN_829 : tag_59; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3918 = _T_5 ? _GEN_830 : tag_60; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3919 = _T_5 ? _GEN_831 : tag_61; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3920 = _T_5 ? _GEN_832 : tag_62; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3921 = _T_5 ? _GEN_833 : tag_63; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3922 = _T_5 ? _GEN_834 : tag_64; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3923 = _T_5 ? _GEN_835 : tag_65; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3924 = _T_5 ? _GEN_836 : tag_66; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3925 = _T_5 ? _GEN_837 : tag_67; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3926 = _T_5 ? _GEN_838 : tag_68; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3927 = _T_5 ? _GEN_839 : tag_69; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3928 = _T_5 ? _GEN_840 : tag_70; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3929 = _T_5 ? _GEN_841 : tag_71; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3930 = _T_5 ? _GEN_842 : tag_72; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3931 = _T_5 ? _GEN_843 : tag_73; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3932 = _T_5 ? _GEN_844 : tag_74; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3933 = _T_5 ? _GEN_845 : tag_75; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3934 = _T_5 ? _GEN_846 : tag_76; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3935 = _T_5 ? _GEN_847 : tag_77; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3936 = _T_5 ? _GEN_848 : tag_78; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3937 = _T_5 ? _GEN_849 : tag_79; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3938 = _T_5 ? _GEN_850 : tag_80; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3939 = _T_5 ? _GEN_851 : tag_81; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3940 = _T_5 ? _GEN_852 : tag_82; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3941 = _T_5 ? _GEN_853 : tag_83; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3942 = _T_5 ? _GEN_854 : tag_84; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3943 = _T_5 ? _GEN_855 : tag_85; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3944 = _T_5 ? _GEN_856 : tag_86; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3945 = _T_5 ? _GEN_857 : tag_87; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3946 = _T_5 ? _GEN_858 : tag_88; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3947 = _T_5 ? _GEN_859 : tag_89; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3948 = _T_5 ? _GEN_860 : tag_90; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3949 = _T_5 ? _GEN_861 : tag_91; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3950 = _T_5 ? _GEN_862 : tag_92; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3951 = _T_5 ? _GEN_863 : tag_93; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3952 = _T_5 ? _GEN_864 : tag_94; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3953 = _T_5 ? _GEN_865 : tag_95; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3954 = _T_5 ? _GEN_866 : tag_96; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3955 = _T_5 ? _GEN_867 : tag_97; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3956 = _T_5 ? _GEN_868 : tag_98; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3957 = _T_5 ? _GEN_869 : tag_99; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3958 = _T_5 ? _GEN_870 : tag_100; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3959 = _T_5 ? _GEN_871 : tag_101; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3960 = _T_5 ? _GEN_872 : tag_102; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3961 = _T_5 ? _GEN_873 : tag_103; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3962 = _T_5 ? _GEN_874 : tag_104; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3963 = _T_5 ? _GEN_875 : tag_105; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3964 = _T_5 ? _GEN_876 : tag_106; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3965 = _T_5 ? _GEN_877 : tag_107; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3966 = _T_5 ? _GEN_878 : tag_108; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3967 = _T_5 ? _GEN_879 : tag_109; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3968 = _T_5 ? _GEN_880 : tag_110; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3969 = _T_5 ? _GEN_881 : tag_111; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3970 = _T_5 ? _GEN_882 : tag_112; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3971 = _T_5 ? _GEN_883 : tag_113; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3972 = _T_5 ? _GEN_884 : tag_114; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3973 = _T_5 ? _GEN_885 : tag_115; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3974 = _T_5 ? _GEN_886 : tag_116; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3975 = _T_5 ? _GEN_887 : tag_117; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3976 = _T_5 ? _GEN_888 : tag_118; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3977 = _T_5 ? _GEN_889 : tag_119; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3978 = _T_5 ? _GEN_890 : tag_120; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3979 = _T_5 ? _GEN_891 : tag_121; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3980 = _T_5 ? _GEN_892 : tag_122; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3981 = _T_5 ? _GEN_893 : tag_123; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3982 = _T_5 ? _GEN_894 : tag_124; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3983 = _T_5 ? _GEN_895 : tag_125; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3984 = _T_5 ? _GEN_896 : tag_126; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3985 = _T_5 ? _GEN_897 : tag_127; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3986 = _T_5 ? _GEN_898 : tag_128; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3987 = _T_5 ? _GEN_899 : tag_129; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3988 = _T_5 ? _GEN_900 : tag_130; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3989 = _T_5 ? _GEN_901 : tag_131; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3990 = _T_5 ? _GEN_902 : tag_132; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3991 = _T_5 ? _GEN_903 : tag_133; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3992 = _T_5 ? _GEN_904 : tag_134; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3993 = _T_5 ? _GEN_905 : tag_135; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3994 = _T_5 ? _GEN_906 : tag_136; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3995 = _T_5 ? _GEN_907 : tag_137; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3996 = _T_5 ? _GEN_908 : tag_138; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3997 = _T_5 ? _GEN_909 : tag_139; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3998 = _T_5 ? _GEN_910 : tag_140; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_3999 = _T_5 ? _GEN_911 : tag_141; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4000 = _T_5 ? _GEN_912 : tag_142; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4001 = _T_5 ? _GEN_913 : tag_143; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4002 = _T_5 ? _GEN_914 : tag_144; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4003 = _T_5 ? _GEN_915 : tag_145; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4004 = _T_5 ? _GEN_916 : tag_146; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4005 = _T_5 ? _GEN_917 : tag_147; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4006 = _T_5 ? _GEN_918 : tag_148; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4007 = _T_5 ? _GEN_919 : tag_149; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4008 = _T_5 ? _GEN_920 : tag_150; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4009 = _T_5 ? _GEN_921 : tag_151; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4010 = _T_5 ? _GEN_922 : tag_152; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4011 = _T_5 ? _GEN_923 : tag_153; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4012 = _T_5 ? _GEN_924 : tag_154; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4013 = _T_5 ? _GEN_925 : tag_155; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4014 = _T_5 ? _GEN_926 : tag_156; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4015 = _T_5 ? _GEN_927 : tag_157; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4016 = _T_5 ? _GEN_928 : tag_158; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4017 = _T_5 ? _GEN_929 : tag_159; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4018 = _T_5 ? _GEN_930 : tag_160; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4019 = _T_5 ? _GEN_931 : tag_161; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4020 = _T_5 ? _GEN_932 : tag_162; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4021 = _T_5 ? _GEN_933 : tag_163; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4022 = _T_5 ? _GEN_934 : tag_164; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4023 = _T_5 ? _GEN_935 : tag_165; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4024 = _T_5 ? _GEN_936 : tag_166; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4025 = _T_5 ? _GEN_937 : tag_167; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4026 = _T_5 ? _GEN_938 : tag_168; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4027 = _T_5 ? _GEN_939 : tag_169; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4028 = _T_5 ? _GEN_940 : tag_170; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4029 = _T_5 ? _GEN_941 : tag_171; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4030 = _T_5 ? _GEN_942 : tag_172; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4031 = _T_5 ? _GEN_943 : tag_173; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4032 = _T_5 ? _GEN_944 : tag_174; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4033 = _T_5 ? _GEN_945 : tag_175; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4034 = _T_5 ? _GEN_946 : tag_176; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4035 = _T_5 ? _GEN_947 : tag_177; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4036 = _T_5 ? _GEN_948 : tag_178; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4037 = _T_5 ? _GEN_949 : tag_179; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4038 = _T_5 ? _GEN_950 : tag_180; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4039 = _T_5 ? _GEN_951 : tag_181; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4040 = _T_5 ? _GEN_952 : tag_182; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4041 = _T_5 ? _GEN_953 : tag_183; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4042 = _T_5 ? _GEN_954 : tag_184; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4043 = _T_5 ? _GEN_955 : tag_185; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4044 = _T_5 ? _GEN_956 : tag_186; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4045 = _T_5 ? _GEN_957 : tag_187; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4046 = _T_5 ? _GEN_958 : tag_188; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4047 = _T_5 ? _GEN_959 : tag_189; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4048 = _T_5 ? _GEN_960 : tag_190; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4049 = _T_5 ? _GEN_961 : tag_191; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4050 = _T_5 ? _GEN_962 : tag_192; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4051 = _T_5 ? _GEN_963 : tag_193; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4052 = _T_5 ? _GEN_964 : tag_194; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4053 = _T_5 ? _GEN_965 : tag_195; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4054 = _T_5 ? _GEN_966 : tag_196; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4055 = _T_5 ? _GEN_967 : tag_197; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4056 = _T_5 ? _GEN_968 : tag_198; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4057 = _T_5 ? _GEN_969 : tag_199; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4058 = _T_5 ? _GEN_970 : tag_200; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4059 = _T_5 ? _GEN_971 : tag_201; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4060 = _T_5 ? _GEN_972 : tag_202; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4061 = _T_5 ? _GEN_973 : tag_203; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4062 = _T_5 ? _GEN_974 : tag_204; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4063 = _T_5 ? _GEN_975 : tag_205; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4064 = _T_5 ? _GEN_976 : tag_206; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4065 = _T_5 ? _GEN_977 : tag_207; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4066 = _T_5 ? _GEN_978 : tag_208; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4067 = _T_5 ? _GEN_979 : tag_209; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4068 = _T_5 ? _GEN_980 : tag_210; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4069 = _T_5 ? _GEN_981 : tag_211; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4070 = _T_5 ? _GEN_982 : tag_212; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4071 = _T_5 ? _GEN_983 : tag_213; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4072 = _T_5 ? _GEN_984 : tag_214; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4073 = _T_5 ? _GEN_985 : tag_215; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4074 = _T_5 ? _GEN_986 : tag_216; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4075 = _T_5 ? _GEN_987 : tag_217; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4076 = _T_5 ? _GEN_988 : tag_218; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4077 = _T_5 ? _GEN_989 : tag_219; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4078 = _T_5 ? _GEN_990 : tag_220; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4079 = _T_5 ? _GEN_991 : tag_221; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4080 = _T_5 ? _GEN_992 : tag_222; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4081 = _T_5 ? _GEN_993 : tag_223; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4082 = _T_5 ? _GEN_994 : tag_224; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4083 = _T_5 ? _GEN_995 : tag_225; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4084 = _T_5 ? _GEN_996 : tag_226; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4085 = _T_5 ? _GEN_997 : tag_227; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4086 = _T_5 ? _GEN_998 : tag_228; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4087 = _T_5 ? _GEN_999 : tag_229; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4088 = _T_5 ? _GEN_1000 : tag_230; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4089 = _T_5 ? _GEN_1001 : tag_231; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4090 = _T_5 ? _GEN_1002 : tag_232; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4091 = _T_5 ? _GEN_1003 : tag_233; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4092 = _T_5 ? _GEN_1004 : tag_234; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4093 = _T_5 ? _GEN_1005 : tag_235; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4094 = _T_5 ? _GEN_1006 : tag_236; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4095 = _T_5 ? _GEN_1007 : tag_237; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4096 = _T_5 ? _GEN_1008 : tag_238; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4097 = _T_5 ? _GEN_1009 : tag_239; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4098 = _T_5 ? _GEN_1010 : tag_240; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4099 = _T_5 ? _GEN_1011 : tag_241; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4100 = _T_5 ? _GEN_1012 : tag_242; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4101 = _T_5 ? _GEN_1013 : tag_243; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4102 = _T_5 ? _GEN_1014 : tag_244; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4103 = _T_5 ? _GEN_1015 : tag_245; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4104 = _T_5 ? _GEN_1016 : tag_246; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4105 = _T_5 ? _GEN_1017 : tag_247; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4106 = _T_5 ? _GEN_1018 : tag_248; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4107 = _T_5 ? _GEN_1019 : tag_249; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4108 = _T_5 ? _GEN_1020 : tag_250; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4109 = _T_5 ? _GEN_1021 : tag_251; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4110 = _T_5 ? _GEN_1022 : tag_252; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4111 = _T_5 ? _GEN_1023 : tag_253; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4112 = _T_5 ? _GEN_1024 : tag_254; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4113 = _T_5 ? _GEN_1025 : tag_255; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [2:0] _GEN_4370 = _T_5 ? 3'h0 : state; // @[Conditional.scala 39:67 Icache.scala 114:25 Icache.scala 26:22]
  wire [2:0] _GEN_4371 = _T_3 ? _GEN_2822 : _GEN_4370; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_4374 = _T_3 ? _GEN_2825 : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_4376 = _T_3 ? _GEN_2827 : _GEN_3599; // @[Conditional.scala 39:67]
  wire  _GEN_4377 = _T_3 ? _GEN_2828 : _GEN_3601; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_4378 = _T_3 ? _GEN_2829 : cache_wdata; // @[Conditional.scala 39:67 Icache.scala 53:28]
  wire  _GEN_4379 = _T_3 ? inst_ready : _GEN_3600; // @[Conditional.scala 39:67 Icache.scala 42:28]
  wire  _GEN_4380 = _T_3 ? valid_0 : _GEN_3602; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4381 = _T_3 ? valid_1 : _GEN_3603; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4382 = _T_3 ? valid_2 : _GEN_3604; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4383 = _T_3 ? valid_3 : _GEN_3605; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4384 = _T_3 ? valid_4 : _GEN_3606; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4385 = _T_3 ? valid_5 : _GEN_3607; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4386 = _T_3 ? valid_6 : _GEN_3608; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4387 = _T_3 ? valid_7 : _GEN_3609; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4388 = _T_3 ? valid_8 : _GEN_3610; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4389 = _T_3 ? valid_9 : _GEN_3611; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4390 = _T_3 ? valid_10 : _GEN_3612; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4391 = _T_3 ? valid_11 : _GEN_3613; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4392 = _T_3 ? valid_12 : _GEN_3614; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4393 = _T_3 ? valid_13 : _GEN_3615; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4394 = _T_3 ? valid_14 : _GEN_3616; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4395 = _T_3 ? valid_15 : _GEN_3617; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4396 = _T_3 ? valid_16 : _GEN_3618; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4397 = _T_3 ? valid_17 : _GEN_3619; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4398 = _T_3 ? valid_18 : _GEN_3620; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4399 = _T_3 ? valid_19 : _GEN_3621; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4400 = _T_3 ? valid_20 : _GEN_3622; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4401 = _T_3 ? valid_21 : _GEN_3623; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4402 = _T_3 ? valid_22 : _GEN_3624; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4403 = _T_3 ? valid_23 : _GEN_3625; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4404 = _T_3 ? valid_24 : _GEN_3626; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4405 = _T_3 ? valid_25 : _GEN_3627; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4406 = _T_3 ? valid_26 : _GEN_3628; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4407 = _T_3 ? valid_27 : _GEN_3629; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4408 = _T_3 ? valid_28 : _GEN_3630; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4409 = _T_3 ? valid_29 : _GEN_3631; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4410 = _T_3 ? valid_30 : _GEN_3632; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4411 = _T_3 ? valid_31 : _GEN_3633; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4412 = _T_3 ? valid_32 : _GEN_3634; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4413 = _T_3 ? valid_33 : _GEN_3635; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4414 = _T_3 ? valid_34 : _GEN_3636; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4415 = _T_3 ? valid_35 : _GEN_3637; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4416 = _T_3 ? valid_36 : _GEN_3638; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4417 = _T_3 ? valid_37 : _GEN_3639; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4418 = _T_3 ? valid_38 : _GEN_3640; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4419 = _T_3 ? valid_39 : _GEN_3641; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4420 = _T_3 ? valid_40 : _GEN_3642; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4421 = _T_3 ? valid_41 : _GEN_3643; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4422 = _T_3 ? valid_42 : _GEN_3644; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4423 = _T_3 ? valid_43 : _GEN_3645; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4424 = _T_3 ? valid_44 : _GEN_3646; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4425 = _T_3 ? valid_45 : _GEN_3647; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4426 = _T_3 ? valid_46 : _GEN_3648; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4427 = _T_3 ? valid_47 : _GEN_3649; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4428 = _T_3 ? valid_48 : _GEN_3650; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4429 = _T_3 ? valid_49 : _GEN_3651; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4430 = _T_3 ? valid_50 : _GEN_3652; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4431 = _T_3 ? valid_51 : _GEN_3653; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4432 = _T_3 ? valid_52 : _GEN_3654; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4433 = _T_3 ? valid_53 : _GEN_3655; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4434 = _T_3 ? valid_54 : _GEN_3656; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4435 = _T_3 ? valid_55 : _GEN_3657; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4436 = _T_3 ? valid_56 : _GEN_3658; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4437 = _T_3 ? valid_57 : _GEN_3659; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4438 = _T_3 ? valid_58 : _GEN_3660; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4439 = _T_3 ? valid_59 : _GEN_3661; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4440 = _T_3 ? valid_60 : _GEN_3662; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4441 = _T_3 ? valid_61 : _GEN_3663; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4442 = _T_3 ? valid_62 : _GEN_3664; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4443 = _T_3 ? valid_63 : _GEN_3665; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4444 = _T_3 ? valid_64 : _GEN_3666; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4445 = _T_3 ? valid_65 : _GEN_3667; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4446 = _T_3 ? valid_66 : _GEN_3668; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4447 = _T_3 ? valid_67 : _GEN_3669; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4448 = _T_3 ? valid_68 : _GEN_3670; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4449 = _T_3 ? valid_69 : _GEN_3671; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4450 = _T_3 ? valid_70 : _GEN_3672; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4451 = _T_3 ? valid_71 : _GEN_3673; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4452 = _T_3 ? valid_72 : _GEN_3674; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4453 = _T_3 ? valid_73 : _GEN_3675; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4454 = _T_3 ? valid_74 : _GEN_3676; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4455 = _T_3 ? valid_75 : _GEN_3677; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4456 = _T_3 ? valid_76 : _GEN_3678; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4457 = _T_3 ? valid_77 : _GEN_3679; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4458 = _T_3 ? valid_78 : _GEN_3680; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4459 = _T_3 ? valid_79 : _GEN_3681; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4460 = _T_3 ? valid_80 : _GEN_3682; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4461 = _T_3 ? valid_81 : _GEN_3683; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4462 = _T_3 ? valid_82 : _GEN_3684; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4463 = _T_3 ? valid_83 : _GEN_3685; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4464 = _T_3 ? valid_84 : _GEN_3686; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4465 = _T_3 ? valid_85 : _GEN_3687; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4466 = _T_3 ? valid_86 : _GEN_3688; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4467 = _T_3 ? valid_87 : _GEN_3689; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4468 = _T_3 ? valid_88 : _GEN_3690; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4469 = _T_3 ? valid_89 : _GEN_3691; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4470 = _T_3 ? valid_90 : _GEN_3692; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4471 = _T_3 ? valid_91 : _GEN_3693; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4472 = _T_3 ? valid_92 : _GEN_3694; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4473 = _T_3 ? valid_93 : _GEN_3695; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4474 = _T_3 ? valid_94 : _GEN_3696; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4475 = _T_3 ? valid_95 : _GEN_3697; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4476 = _T_3 ? valid_96 : _GEN_3698; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4477 = _T_3 ? valid_97 : _GEN_3699; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4478 = _T_3 ? valid_98 : _GEN_3700; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4479 = _T_3 ? valid_99 : _GEN_3701; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4480 = _T_3 ? valid_100 : _GEN_3702; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4481 = _T_3 ? valid_101 : _GEN_3703; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4482 = _T_3 ? valid_102 : _GEN_3704; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4483 = _T_3 ? valid_103 : _GEN_3705; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4484 = _T_3 ? valid_104 : _GEN_3706; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4485 = _T_3 ? valid_105 : _GEN_3707; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4486 = _T_3 ? valid_106 : _GEN_3708; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4487 = _T_3 ? valid_107 : _GEN_3709; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4488 = _T_3 ? valid_108 : _GEN_3710; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4489 = _T_3 ? valid_109 : _GEN_3711; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4490 = _T_3 ? valid_110 : _GEN_3712; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4491 = _T_3 ? valid_111 : _GEN_3713; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4492 = _T_3 ? valid_112 : _GEN_3714; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4493 = _T_3 ? valid_113 : _GEN_3715; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4494 = _T_3 ? valid_114 : _GEN_3716; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4495 = _T_3 ? valid_115 : _GEN_3717; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4496 = _T_3 ? valid_116 : _GEN_3718; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4497 = _T_3 ? valid_117 : _GEN_3719; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4498 = _T_3 ? valid_118 : _GEN_3720; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4499 = _T_3 ? valid_119 : _GEN_3721; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4500 = _T_3 ? valid_120 : _GEN_3722; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4501 = _T_3 ? valid_121 : _GEN_3723; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4502 = _T_3 ? valid_122 : _GEN_3724; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4503 = _T_3 ? valid_123 : _GEN_3725; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4504 = _T_3 ? valid_124 : _GEN_3726; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4505 = _T_3 ? valid_125 : _GEN_3727; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4506 = _T_3 ? valid_126 : _GEN_3728; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4507 = _T_3 ? valid_127 : _GEN_3729; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4508 = _T_3 ? valid_128 : _GEN_3730; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4509 = _T_3 ? valid_129 : _GEN_3731; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4510 = _T_3 ? valid_130 : _GEN_3732; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4511 = _T_3 ? valid_131 : _GEN_3733; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4512 = _T_3 ? valid_132 : _GEN_3734; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4513 = _T_3 ? valid_133 : _GEN_3735; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4514 = _T_3 ? valid_134 : _GEN_3736; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4515 = _T_3 ? valid_135 : _GEN_3737; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4516 = _T_3 ? valid_136 : _GEN_3738; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4517 = _T_3 ? valid_137 : _GEN_3739; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4518 = _T_3 ? valid_138 : _GEN_3740; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4519 = _T_3 ? valid_139 : _GEN_3741; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4520 = _T_3 ? valid_140 : _GEN_3742; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4521 = _T_3 ? valid_141 : _GEN_3743; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4522 = _T_3 ? valid_142 : _GEN_3744; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4523 = _T_3 ? valid_143 : _GEN_3745; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4524 = _T_3 ? valid_144 : _GEN_3746; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4525 = _T_3 ? valid_145 : _GEN_3747; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4526 = _T_3 ? valid_146 : _GEN_3748; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4527 = _T_3 ? valid_147 : _GEN_3749; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4528 = _T_3 ? valid_148 : _GEN_3750; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4529 = _T_3 ? valid_149 : _GEN_3751; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4530 = _T_3 ? valid_150 : _GEN_3752; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4531 = _T_3 ? valid_151 : _GEN_3753; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4532 = _T_3 ? valid_152 : _GEN_3754; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4533 = _T_3 ? valid_153 : _GEN_3755; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4534 = _T_3 ? valid_154 : _GEN_3756; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4535 = _T_3 ? valid_155 : _GEN_3757; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4536 = _T_3 ? valid_156 : _GEN_3758; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4537 = _T_3 ? valid_157 : _GEN_3759; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4538 = _T_3 ? valid_158 : _GEN_3760; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4539 = _T_3 ? valid_159 : _GEN_3761; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4540 = _T_3 ? valid_160 : _GEN_3762; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4541 = _T_3 ? valid_161 : _GEN_3763; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4542 = _T_3 ? valid_162 : _GEN_3764; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4543 = _T_3 ? valid_163 : _GEN_3765; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4544 = _T_3 ? valid_164 : _GEN_3766; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4545 = _T_3 ? valid_165 : _GEN_3767; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4546 = _T_3 ? valid_166 : _GEN_3768; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4547 = _T_3 ? valid_167 : _GEN_3769; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4548 = _T_3 ? valid_168 : _GEN_3770; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4549 = _T_3 ? valid_169 : _GEN_3771; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4550 = _T_3 ? valid_170 : _GEN_3772; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4551 = _T_3 ? valid_171 : _GEN_3773; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4552 = _T_3 ? valid_172 : _GEN_3774; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4553 = _T_3 ? valid_173 : _GEN_3775; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4554 = _T_3 ? valid_174 : _GEN_3776; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4555 = _T_3 ? valid_175 : _GEN_3777; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4556 = _T_3 ? valid_176 : _GEN_3778; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4557 = _T_3 ? valid_177 : _GEN_3779; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4558 = _T_3 ? valid_178 : _GEN_3780; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4559 = _T_3 ? valid_179 : _GEN_3781; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4560 = _T_3 ? valid_180 : _GEN_3782; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4561 = _T_3 ? valid_181 : _GEN_3783; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4562 = _T_3 ? valid_182 : _GEN_3784; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4563 = _T_3 ? valid_183 : _GEN_3785; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4564 = _T_3 ? valid_184 : _GEN_3786; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4565 = _T_3 ? valid_185 : _GEN_3787; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4566 = _T_3 ? valid_186 : _GEN_3788; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4567 = _T_3 ? valid_187 : _GEN_3789; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4568 = _T_3 ? valid_188 : _GEN_3790; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4569 = _T_3 ? valid_189 : _GEN_3791; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4570 = _T_3 ? valid_190 : _GEN_3792; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4571 = _T_3 ? valid_191 : _GEN_3793; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4572 = _T_3 ? valid_192 : _GEN_3794; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4573 = _T_3 ? valid_193 : _GEN_3795; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4574 = _T_3 ? valid_194 : _GEN_3796; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4575 = _T_3 ? valid_195 : _GEN_3797; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4576 = _T_3 ? valid_196 : _GEN_3798; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4577 = _T_3 ? valid_197 : _GEN_3799; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4578 = _T_3 ? valid_198 : _GEN_3800; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4579 = _T_3 ? valid_199 : _GEN_3801; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4580 = _T_3 ? valid_200 : _GEN_3802; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4581 = _T_3 ? valid_201 : _GEN_3803; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4582 = _T_3 ? valid_202 : _GEN_3804; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4583 = _T_3 ? valid_203 : _GEN_3805; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4584 = _T_3 ? valid_204 : _GEN_3806; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4585 = _T_3 ? valid_205 : _GEN_3807; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4586 = _T_3 ? valid_206 : _GEN_3808; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4587 = _T_3 ? valid_207 : _GEN_3809; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4588 = _T_3 ? valid_208 : _GEN_3810; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4589 = _T_3 ? valid_209 : _GEN_3811; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4590 = _T_3 ? valid_210 : _GEN_3812; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4591 = _T_3 ? valid_211 : _GEN_3813; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4592 = _T_3 ? valid_212 : _GEN_3814; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4593 = _T_3 ? valid_213 : _GEN_3815; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4594 = _T_3 ? valid_214 : _GEN_3816; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4595 = _T_3 ? valid_215 : _GEN_3817; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4596 = _T_3 ? valid_216 : _GEN_3818; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4597 = _T_3 ? valid_217 : _GEN_3819; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4598 = _T_3 ? valid_218 : _GEN_3820; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4599 = _T_3 ? valid_219 : _GEN_3821; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4600 = _T_3 ? valid_220 : _GEN_3822; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4601 = _T_3 ? valid_221 : _GEN_3823; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4602 = _T_3 ? valid_222 : _GEN_3824; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4603 = _T_3 ? valid_223 : _GEN_3825; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4604 = _T_3 ? valid_224 : _GEN_3826; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4605 = _T_3 ? valid_225 : _GEN_3827; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4606 = _T_3 ? valid_226 : _GEN_3828; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4607 = _T_3 ? valid_227 : _GEN_3829; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4608 = _T_3 ? valid_228 : _GEN_3830; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4609 = _T_3 ? valid_229 : _GEN_3831; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4610 = _T_3 ? valid_230 : _GEN_3832; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4611 = _T_3 ? valid_231 : _GEN_3833; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4612 = _T_3 ? valid_232 : _GEN_3834; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4613 = _T_3 ? valid_233 : _GEN_3835; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4614 = _T_3 ? valid_234 : _GEN_3836; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4615 = _T_3 ? valid_235 : _GEN_3837; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4616 = _T_3 ? valid_236 : _GEN_3838; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4617 = _T_3 ? valid_237 : _GEN_3839; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4618 = _T_3 ? valid_238 : _GEN_3840; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4619 = _T_3 ? valid_239 : _GEN_3841; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4620 = _T_3 ? valid_240 : _GEN_3842; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4621 = _T_3 ? valid_241 : _GEN_3843; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4622 = _T_3 ? valid_242 : _GEN_3844; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4623 = _T_3 ? valid_243 : _GEN_3845; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4624 = _T_3 ? valid_244 : _GEN_3846; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4625 = _T_3 ? valid_245 : _GEN_3847; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4626 = _T_3 ? valid_246 : _GEN_3848; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4627 = _T_3 ? valid_247 : _GEN_3849; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4628 = _T_3 ? valid_248 : _GEN_3850; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4629 = _T_3 ? valid_249 : _GEN_3851; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4630 = _T_3 ? valid_250 : _GEN_3852; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4631 = _T_3 ? valid_251 : _GEN_3853; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4632 = _T_3 ? valid_252 : _GEN_3854; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4633 = _T_3 ? valid_253 : _GEN_3855; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4634 = _T_3 ? valid_254 : _GEN_3856; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire  _GEN_4635 = _T_3 ? valid_255 : _GEN_3857; // @[Conditional.scala 39:67 Icache.scala 18:24]
  wire [19:0] _GEN_4636 = _T_3 ? tag_0 : _GEN_3858; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4637 = _T_3 ? tag_1 : _GEN_3859; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4638 = _T_3 ? tag_2 : _GEN_3860; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4639 = _T_3 ? tag_3 : _GEN_3861; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4640 = _T_3 ? tag_4 : _GEN_3862; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4641 = _T_3 ? tag_5 : _GEN_3863; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4642 = _T_3 ? tag_6 : _GEN_3864; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4643 = _T_3 ? tag_7 : _GEN_3865; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4644 = _T_3 ? tag_8 : _GEN_3866; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4645 = _T_3 ? tag_9 : _GEN_3867; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4646 = _T_3 ? tag_10 : _GEN_3868; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4647 = _T_3 ? tag_11 : _GEN_3869; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4648 = _T_3 ? tag_12 : _GEN_3870; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4649 = _T_3 ? tag_13 : _GEN_3871; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4650 = _T_3 ? tag_14 : _GEN_3872; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4651 = _T_3 ? tag_15 : _GEN_3873; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4652 = _T_3 ? tag_16 : _GEN_3874; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4653 = _T_3 ? tag_17 : _GEN_3875; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4654 = _T_3 ? tag_18 : _GEN_3876; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4655 = _T_3 ? tag_19 : _GEN_3877; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4656 = _T_3 ? tag_20 : _GEN_3878; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4657 = _T_3 ? tag_21 : _GEN_3879; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4658 = _T_3 ? tag_22 : _GEN_3880; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4659 = _T_3 ? tag_23 : _GEN_3881; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4660 = _T_3 ? tag_24 : _GEN_3882; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4661 = _T_3 ? tag_25 : _GEN_3883; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4662 = _T_3 ? tag_26 : _GEN_3884; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4663 = _T_3 ? tag_27 : _GEN_3885; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4664 = _T_3 ? tag_28 : _GEN_3886; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4665 = _T_3 ? tag_29 : _GEN_3887; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4666 = _T_3 ? tag_30 : _GEN_3888; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4667 = _T_3 ? tag_31 : _GEN_3889; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4668 = _T_3 ? tag_32 : _GEN_3890; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4669 = _T_3 ? tag_33 : _GEN_3891; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4670 = _T_3 ? tag_34 : _GEN_3892; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4671 = _T_3 ? tag_35 : _GEN_3893; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4672 = _T_3 ? tag_36 : _GEN_3894; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4673 = _T_3 ? tag_37 : _GEN_3895; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4674 = _T_3 ? tag_38 : _GEN_3896; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4675 = _T_3 ? tag_39 : _GEN_3897; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4676 = _T_3 ? tag_40 : _GEN_3898; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4677 = _T_3 ? tag_41 : _GEN_3899; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4678 = _T_3 ? tag_42 : _GEN_3900; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4679 = _T_3 ? tag_43 : _GEN_3901; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4680 = _T_3 ? tag_44 : _GEN_3902; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4681 = _T_3 ? tag_45 : _GEN_3903; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4682 = _T_3 ? tag_46 : _GEN_3904; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4683 = _T_3 ? tag_47 : _GEN_3905; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4684 = _T_3 ? tag_48 : _GEN_3906; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4685 = _T_3 ? tag_49 : _GEN_3907; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4686 = _T_3 ? tag_50 : _GEN_3908; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4687 = _T_3 ? tag_51 : _GEN_3909; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4688 = _T_3 ? tag_52 : _GEN_3910; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4689 = _T_3 ? tag_53 : _GEN_3911; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4690 = _T_3 ? tag_54 : _GEN_3912; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4691 = _T_3 ? tag_55 : _GEN_3913; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4692 = _T_3 ? tag_56 : _GEN_3914; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4693 = _T_3 ? tag_57 : _GEN_3915; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4694 = _T_3 ? tag_58 : _GEN_3916; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4695 = _T_3 ? tag_59 : _GEN_3917; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4696 = _T_3 ? tag_60 : _GEN_3918; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4697 = _T_3 ? tag_61 : _GEN_3919; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4698 = _T_3 ? tag_62 : _GEN_3920; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4699 = _T_3 ? tag_63 : _GEN_3921; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4700 = _T_3 ? tag_64 : _GEN_3922; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4701 = _T_3 ? tag_65 : _GEN_3923; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4702 = _T_3 ? tag_66 : _GEN_3924; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4703 = _T_3 ? tag_67 : _GEN_3925; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4704 = _T_3 ? tag_68 : _GEN_3926; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4705 = _T_3 ? tag_69 : _GEN_3927; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4706 = _T_3 ? tag_70 : _GEN_3928; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4707 = _T_3 ? tag_71 : _GEN_3929; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4708 = _T_3 ? tag_72 : _GEN_3930; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4709 = _T_3 ? tag_73 : _GEN_3931; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4710 = _T_3 ? tag_74 : _GEN_3932; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4711 = _T_3 ? tag_75 : _GEN_3933; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4712 = _T_3 ? tag_76 : _GEN_3934; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4713 = _T_3 ? tag_77 : _GEN_3935; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4714 = _T_3 ? tag_78 : _GEN_3936; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4715 = _T_3 ? tag_79 : _GEN_3937; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4716 = _T_3 ? tag_80 : _GEN_3938; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4717 = _T_3 ? tag_81 : _GEN_3939; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4718 = _T_3 ? tag_82 : _GEN_3940; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4719 = _T_3 ? tag_83 : _GEN_3941; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4720 = _T_3 ? tag_84 : _GEN_3942; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4721 = _T_3 ? tag_85 : _GEN_3943; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4722 = _T_3 ? tag_86 : _GEN_3944; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4723 = _T_3 ? tag_87 : _GEN_3945; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4724 = _T_3 ? tag_88 : _GEN_3946; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4725 = _T_3 ? tag_89 : _GEN_3947; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4726 = _T_3 ? tag_90 : _GEN_3948; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4727 = _T_3 ? tag_91 : _GEN_3949; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4728 = _T_3 ? tag_92 : _GEN_3950; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4729 = _T_3 ? tag_93 : _GEN_3951; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4730 = _T_3 ? tag_94 : _GEN_3952; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4731 = _T_3 ? tag_95 : _GEN_3953; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4732 = _T_3 ? tag_96 : _GEN_3954; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4733 = _T_3 ? tag_97 : _GEN_3955; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4734 = _T_3 ? tag_98 : _GEN_3956; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4735 = _T_3 ? tag_99 : _GEN_3957; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4736 = _T_3 ? tag_100 : _GEN_3958; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4737 = _T_3 ? tag_101 : _GEN_3959; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4738 = _T_3 ? tag_102 : _GEN_3960; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4739 = _T_3 ? tag_103 : _GEN_3961; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4740 = _T_3 ? tag_104 : _GEN_3962; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4741 = _T_3 ? tag_105 : _GEN_3963; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4742 = _T_3 ? tag_106 : _GEN_3964; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4743 = _T_3 ? tag_107 : _GEN_3965; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4744 = _T_3 ? tag_108 : _GEN_3966; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4745 = _T_3 ? tag_109 : _GEN_3967; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4746 = _T_3 ? tag_110 : _GEN_3968; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4747 = _T_3 ? tag_111 : _GEN_3969; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4748 = _T_3 ? tag_112 : _GEN_3970; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4749 = _T_3 ? tag_113 : _GEN_3971; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4750 = _T_3 ? tag_114 : _GEN_3972; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4751 = _T_3 ? tag_115 : _GEN_3973; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4752 = _T_3 ? tag_116 : _GEN_3974; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4753 = _T_3 ? tag_117 : _GEN_3975; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4754 = _T_3 ? tag_118 : _GEN_3976; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4755 = _T_3 ? tag_119 : _GEN_3977; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4756 = _T_3 ? tag_120 : _GEN_3978; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4757 = _T_3 ? tag_121 : _GEN_3979; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4758 = _T_3 ? tag_122 : _GEN_3980; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4759 = _T_3 ? tag_123 : _GEN_3981; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4760 = _T_3 ? tag_124 : _GEN_3982; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4761 = _T_3 ? tag_125 : _GEN_3983; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4762 = _T_3 ? tag_126 : _GEN_3984; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4763 = _T_3 ? tag_127 : _GEN_3985; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4764 = _T_3 ? tag_128 : _GEN_3986; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4765 = _T_3 ? tag_129 : _GEN_3987; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4766 = _T_3 ? tag_130 : _GEN_3988; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4767 = _T_3 ? tag_131 : _GEN_3989; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4768 = _T_3 ? tag_132 : _GEN_3990; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4769 = _T_3 ? tag_133 : _GEN_3991; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4770 = _T_3 ? tag_134 : _GEN_3992; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4771 = _T_3 ? tag_135 : _GEN_3993; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4772 = _T_3 ? tag_136 : _GEN_3994; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4773 = _T_3 ? tag_137 : _GEN_3995; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4774 = _T_3 ? tag_138 : _GEN_3996; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4775 = _T_3 ? tag_139 : _GEN_3997; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4776 = _T_3 ? tag_140 : _GEN_3998; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4777 = _T_3 ? tag_141 : _GEN_3999; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4778 = _T_3 ? tag_142 : _GEN_4000; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4779 = _T_3 ? tag_143 : _GEN_4001; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4780 = _T_3 ? tag_144 : _GEN_4002; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4781 = _T_3 ? tag_145 : _GEN_4003; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4782 = _T_3 ? tag_146 : _GEN_4004; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4783 = _T_3 ? tag_147 : _GEN_4005; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4784 = _T_3 ? tag_148 : _GEN_4006; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4785 = _T_3 ? tag_149 : _GEN_4007; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4786 = _T_3 ? tag_150 : _GEN_4008; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4787 = _T_3 ? tag_151 : _GEN_4009; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4788 = _T_3 ? tag_152 : _GEN_4010; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4789 = _T_3 ? tag_153 : _GEN_4011; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4790 = _T_3 ? tag_154 : _GEN_4012; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4791 = _T_3 ? tag_155 : _GEN_4013; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4792 = _T_3 ? tag_156 : _GEN_4014; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4793 = _T_3 ? tag_157 : _GEN_4015; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4794 = _T_3 ? tag_158 : _GEN_4016; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4795 = _T_3 ? tag_159 : _GEN_4017; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4796 = _T_3 ? tag_160 : _GEN_4018; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4797 = _T_3 ? tag_161 : _GEN_4019; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4798 = _T_3 ? tag_162 : _GEN_4020; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4799 = _T_3 ? tag_163 : _GEN_4021; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4800 = _T_3 ? tag_164 : _GEN_4022; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4801 = _T_3 ? tag_165 : _GEN_4023; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4802 = _T_3 ? tag_166 : _GEN_4024; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4803 = _T_3 ? tag_167 : _GEN_4025; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4804 = _T_3 ? tag_168 : _GEN_4026; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4805 = _T_3 ? tag_169 : _GEN_4027; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4806 = _T_3 ? tag_170 : _GEN_4028; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4807 = _T_3 ? tag_171 : _GEN_4029; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4808 = _T_3 ? tag_172 : _GEN_4030; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4809 = _T_3 ? tag_173 : _GEN_4031; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4810 = _T_3 ? tag_174 : _GEN_4032; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4811 = _T_3 ? tag_175 : _GEN_4033; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4812 = _T_3 ? tag_176 : _GEN_4034; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4813 = _T_3 ? tag_177 : _GEN_4035; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4814 = _T_3 ? tag_178 : _GEN_4036; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4815 = _T_3 ? tag_179 : _GEN_4037; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4816 = _T_3 ? tag_180 : _GEN_4038; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4817 = _T_3 ? tag_181 : _GEN_4039; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4818 = _T_3 ? tag_182 : _GEN_4040; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4819 = _T_3 ? tag_183 : _GEN_4041; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4820 = _T_3 ? tag_184 : _GEN_4042; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4821 = _T_3 ? tag_185 : _GEN_4043; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4822 = _T_3 ? tag_186 : _GEN_4044; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4823 = _T_3 ? tag_187 : _GEN_4045; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4824 = _T_3 ? tag_188 : _GEN_4046; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4825 = _T_3 ? tag_189 : _GEN_4047; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4826 = _T_3 ? tag_190 : _GEN_4048; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4827 = _T_3 ? tag_191 : _GEN_4049; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4828 = _T_3 ? tag_192 : _GEN_4050; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4829 = _T_3 ? tag_193 : _GEN_4051; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4830 = _T_3 ? tag_194 : _GEN_4052; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4831 = _T_3 ? tag_195 : _GEN_4053; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4832 = _T_3 ? tag_196 : _GEN_4054; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4833 = _T_3 ? tag_197 : _GEN_4055; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4834 = _T_3 ? tag_198 : _GEN_4056; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4835 = _T_3 ? tag_199 : _GEN_4057; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4836 = _T_3 ? tag_200 : _GEN_4058; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4837 = _T_3 ? tag_201 : _GEN_4059; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4838 = _T_3 ? tag_202 : _GEN_4060; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4839 = _T_3 ? tag_203 : _GEN_4061; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4840 = _T_3 ? tag_204 : _GEN_4062; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4841 = _T_3 ? tag_205 : _GEN_4063; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4842 = _T_3 ? tag_206 : _GEN_4064; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4843 = _T_3 ? tag_207 : _GEN_4065; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4844 = _T_3 ? tag_208 : _GEN_4066; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4845 = _T_3 ? tag_209 : _GEN_4067; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4846 = _T_3 ? tag_210 : _GEN_4068; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4847 = _T_3 ? tag_211 : _GEN_4069; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4848 = _T_3 ? tag_212 : _GEN_4070; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4849 = _T_3 ? tag_213 : _GEN_4071; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4850 = _T_3 ? tag_214 : _GEN_4072; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4851 = _T_3 ? tag_215 : _GEN_4073; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4852 = _T_3 ? tag_216 : _GEN_4074; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4853 = _T_3 ? tag_217 : _GEN_4075; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4854 = _T_3 ? tag_218 : _GEN_4076; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4855 = _T_3 ? tag_219 : _GEN_4077; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4856 = _T_3 ? tag_220 : _GEN_4078; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4857 = _T_3 ? tag_221 : _GEN_4079; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4858 = _T_3 ? tag_222 : _GEN_4080; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4859 = _T_3 ? tag_223 : _GEN_4081; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4860 = _T_3 ? tag_224 : _GEN_4082; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4861 = _T_3 ? tag_225 : _GEN_4083; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4862 = _T_3 ? tag_226 : _GEN_4084; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4863 = _T_3 ? tag_227 : _GEN_4085; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4864 = _T_3 ? tag_228 : _GEN_4086; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4865 = _T_3 ? tag_229 : _GEN_4087; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4866 = _T_3 ? tag_230 : _GEN_4088; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4867 = _T_3 ? tag_231 : _GEN_4089; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4868 = _T_3 ? tag_232 : _GEN_4090; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4869 = _T_3 ? tag_233 : _GEN_4091; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4870 = _T_3 ? tag_234 : _GEN_4092; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4871 = _T_3 ? tag_235 : _GEN_4093; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4872 = _T_3 ? tag_236 : _GEN_4094; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4873 = _T_3 ? tag_237 : _GEN_4095; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4874 = _T_3 ? tag_238 : _GEN_4096; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4875 = _T_3 ? tag_239 : _GEN_4097; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4876 = _T_3 ? tag_240 : _GEN_4098; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4877 = _T_3 ? tag_241 : _GEN_4099; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4878 = _T_3 ? tag_242 : _GEN_4100; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4879 = _T_3 ? tag_243 : _GEN_4101; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4880 = _T_3 ? tag_244 : _GEN_4102; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4881 = _T_3 ? tag_245 : _GEN_4103; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4882 = _T_3 ? tag_246 : _GEN_4104; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4883 = _T_3 ? tag_247 : _GEN_4105; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4884 = _T_3 ? tag_248 : _GEN_4106; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4885 = _T_3 ? tag_249 : _GEN_4107; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4886 = _T_3 ? tag_250 : _GEN_4108; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4887 = _T_3 ? tag_251 : _GEN_4109; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4888 = _T_3 ? tag_252 : _GEN_4110; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4889 = _T_3 ? tag_253 : _GEN_4111; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4890 = _T_3 ? tag_254 : _GEN_4112; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_4891 = _T_3 ? tag_255 : _GEN_4113; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_5918 = _T_2 ? 1'h0 : _T_3 & _GEN_2830; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_5920 = _T_2 ? 32'h0 : _GEN_4374; // @[Conditional.scala 39:67]
  wire  _GEN_6695 = _T_1 ? 1'h0 : _GEN_5918; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_6697 = _T_1 ? 32'h0 : _GEN_5920; // @[Conditional.scala 39:67]
  S011HD1P_X32Y2D128 req ( // @[Icache.scala 126:19]
    .Q(req_Q),
    .CLK(req_CLK),
    .CEN(req_CEN),
    .WEN(req_WEN),
    .A(req_A),
    .D(req_D)
  );
  assign io_imem_inst_ready = inst_ready; // @[Icache.scala 123:19]
  assign io_imem_inst_read = 2'h3 == req_offset[3:2] ? cache_data_out[127:96] : _inst_read_T_8; // @[Mux.scala 80:57]
  assign io_out_inst_valid = _T ? 1'h0 : _GEN_6695; // @[Conditional.scala 40:58]
  assign io_out_inst_addr = _T ? 32'h0 : _GEN_6697; // @[Conditional.scala 40:58]
  assign req_CLK = clock; // @[Icache.scala 127:14]
  assign req_CEN = 1'h1; // @[Icache.scala 128:14]
  assign req_WEN = cache_wen; // @[Icache.scala 129:14]
  assign req_A = io_imem_inst_addr[11:4]; // @[Icache.scala 29:30]
  assign req_D = cache_wdata; // @[Icache.scala 131:14]
  always @(posedge clock) begin
    if (reset) begin // @[Icache.scala 17:24]
      tag_0 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_0 <= _GEN_2309;
        end else begin
          tag_0 <= _GEN_4636;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_1 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_1 <= _GEN_2310;
        end else begin
          tag_1 <= _GEN_4637;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_2 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_2 <= _GEN_2311;
        end else begin
          tag_2 <= _GEN_4638;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_3 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_3 <= _GEN_2312;
        end else begin
          tag_3 <= _GEN_4639;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_4 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_4 <= _GEN_2313;
        end else begin
          tag_4 <= _GEN_4640;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_5 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_5 <= _GEN_2314;
        end else begin
          tag_5 <= _GEN_4641;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_6 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_6 <= _GEN_2315;
        end else begin
          tag_6 <= _GEN_4642;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_7 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_7 <= _GEN_2316;
        end else begin
          tag_7 <= _GEN_4643;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_8 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_8 <= _GEN_2317;
        end else begin
          tag_8 <= _GEN_4644;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_9 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_9 <= _GEN_2318;
        end else begin
          tag_9 <= _GEN_4645;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_10 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_10 <= _GEN_2319;
        end else begin
          tag_10 <= _GEN_4646;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_11 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_11 <= _GEN_2320;
        end else begin
          tag_11 <= _GEN_4647;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_12 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_12 <= _GEN_2321;
        end else begin
          tag_12 <= _GEN_4648;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_13 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_13 <= _GEN_2322;
        end else begin
          tag_13 <= _GEN_4649;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_14 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_14 <= _GEN_2323;
        end else begin
          tag_14 <= _GEN_4650;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_15 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_15 <= _GEN_2324;
        end else begin
          tag_15 <= _GEN_4651;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_16 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_16 <= _GEN_2325;
        end else begin
          tag_16 <= _GEN_4652;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_17 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_17 <= _GEN_2326;
        end else begin
          tag_17 <= _GEN_4653;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_18 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_18 <= _GEN_2327;
        end else begin
          tag_18 <= _GEN_4654;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_19 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_19 <= _GEN_2328;
        end else begin
          tag_19 <= _GEN_4655;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_20 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_20 <= _GEN_2329;
        end else begin
          tag_20 <= _GEN_4656;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_21 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_21 <= _GEN_2330;
        end else begin
          tag_21 <= _GEN_4657;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_22 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_22 <= _GEN_2331;
        end else begin
          tag_22 <= _GEN_4658;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_23 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_23 <= _GEN_2332;
        end else begin
          tag_23 <= _GEN_4659;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_24 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_24 <= _GEN_2333;
        end else begin
          tag_24 <= _GEN_4660;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_25 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_25 <= _GEN_2334;
        end else begin
          tag_25 <= _GEN_4661;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_26 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_26 <= _GEN_2335;
        end else begin
          tag_26 <= _GEN_4662;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_27 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_27 <= _GEN_2336;
        end else begin
          tag_27 <= _GEN_4663;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_28 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_28 <= _GEN_2337;
        end else begin
          tag_28 <= _GEN_4664;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_29 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_29 <= _GEN_2338;
        end else begin
          tag_29 <= _GEN_4665;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_30 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_30 <= _GEN_2339;
        end else begin
          tag_30 <= _GEN_4666;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_31 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_31 <= _GEN_2340;
        end else begin
          tag_31 <= _GEN_4667;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_32 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_32 <= _GEN_2341;
        end else begin
          tag_32 <= _GEN_4668;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_33 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_33 <= _GEN_2342;
        end else begin
          tag_33 <= _GEN_4669;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_34 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_34 <= _GEN_2343;
        end else begin
          tag_34 <= _GEN_4670;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_35 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_35 <= _GEN_2344;
        end else begin
          tag_35 <= _GEN_4671;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_36 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_36 <= _GEN_2345;
        end else begin
          tag_36 <= _GEN_4672;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_37 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_37 <= _GEN_2346;
        end else begin
          tag_37 <= _GEN_4673;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_38 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_38 <= _GEN_2347;
        end else begin
          tag_38 <= _GEN_4674;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_39 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_39 <= _GEN_2348;
        end else begin
          tag_39 <= _GEN_4675;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_40 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_40 <= _GEN_2349;
        end else begin
          tag_40 <= _GEN_4676;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_41 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_41 <= _GEN_2350;
        end else begin
          tag_41 <= _GEN_4677;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_42 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_42 <= _GEN_2351;
        end else begin
          tag_42 <= _GEN_4678;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_43 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_43 <= _GEN_2352;
        end else begin
          tag_43 <= _GEN_4679;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_44 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_44 <= _GEN_2353;
        end else begin
          tag_44 <= _GEN_4680;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_45 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_45 <= _GEN_2354;
        end else begin
          tag_45 <= _GEN_4681;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_46 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_46 <= _GEN_2355;
        end else begin
          tag_46 <= _GEN_4682;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_47 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_47 <= _GEN_2356;
        end else begin
          tag_47 <= _GEN_4683;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_48 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_48 <= _GEN_2357;
        end else begin
          tag_48 <= _GEN_4684;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_49 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_49 <= _GEN_2358;
        end else begin
          tag_49 <= _GEN_4685;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_50 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_50 <= _GEN_2359;
        end else begin
          tag_50 <= _GEN_4686;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_51 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_51 <= _GEN_2360;
        end else begin
          tag_51 <= _GEN_4687;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_52 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_52 <= _GEN_2361;
        end else begin
          tag_52 <= _GEN_4688;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_53 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_53 <= _GEN_2362;
        end else begin
          tag_53 <= _GEN_4689;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_54 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_54 <= _GEN_2363;
        end else begin
          tag_54 <= _GEN_4690;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_55 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_55 <= _GEN_2364;
        end else begin
          tag_55 <= _GEN_4691;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_56 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_56 <= _GEN_2365;
        end else begin
          tag_56 <= _GEN_4692;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_57 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_57 <= _GEN_2366;
        end else begin
          tag_57 <= _GEN_4693;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_58 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_58 <= _GEN_2367;
        end else begin
          tag_58 <= _GEN_4694;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_59 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_59 <= _GEN_2368;
        end else begin
          tag_59 <= _GEN_4695;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_60 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_60 <= _GEN_2369;
        end else begin
          tag_60 <= _GEN_4696;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_61 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_61 <= _GEN_2370;
        end else begin
          tag_61 <= _GEN_4697;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_62 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_62 <= _GEN_2371;
        end else begin
          tag_62 <= _GEN_4698;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_63 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_63 <= _GEN_2372;
        end else begin
          tag_63 <= _GEN_4699;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_64 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_64 <= _GEN_2373;
        end else begin
          tag_64 <= _GEN_4700;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_65 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_65 <= _GEN_2374;
        end else begin
          tag_65 <= _GEN_4701;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_66 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_66 <= _GEN_2375;
        end else begin
          tag_66 <= _GEN_4702;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_67 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_67 <= _GEN_2376;
        end else begin
          tag_67 <= _GEN_4703;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_68 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_68 <= _GEN_2377;
        end else begin
          tag_68 <= _GEN_4704;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_69 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_69 <= _GEN_2378;
        end else begin
          tag_69 <= _GEN_4705;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_70 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_70 <= _GEN_2379;
        end else begin
          tag_70 <= _GEN_4706;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_71 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_71 <= _GEN_2380;
        end else begin
          tag_71 <= _GEN_4707;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_72 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_72 <= _GEN_2381;
        end else begin
          tag_72 <= _GEN_4708;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_73 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_73 <= _GEN_2382;
        end else begin
          tag_73 <= _GEN_4709;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_74 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_74 <= _GEN_2383;
        end else begin
          tag_74 <= _GEN_4710;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_75 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_75 <= _GEN_2384;
        end else begin
          tag_75 <= _GEN_4711;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_76 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_76 <= _GEN_2385;
        end else begin
          tag_76 <= _GEN_4712;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_77 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_77 <= _GEN_2386;
        end else begin
          tag_77 <= _GEN_4713;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_78 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_78 <= _GEN_2387;
        end else begin
          tag_78 <= _GEN_4714;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_79 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_79 <= _GEN_2388;
        end else begin
          tag_79 <= _GEN_4715;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_80 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_80 <= _GEN_2389;
        end else begin
          tag_80 <= _GEN_4716;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_81 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_81 <= _GEN_2390;
        end else begin
          tag_81 <= _GEN_4717;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_82 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_82 <= _GEN_2391;
        end else begin
          tag_82 <= _GEN_4718;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_83 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_83 <= _GEN_2392;
        end else begin
          tag_83 <= _GEN_4719;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_84 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_84 <= _GEN_2393;
        end else begin
          tag_84 <= _GEN_4720;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_85 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_85 <= _GEN_2394;
        end else begin
          tag_85 <= _GEN_4721;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_86 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_86 <= _GEN_2395;
        end else begin
          tag_86 <= _GEN_4722;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_87 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_87 <= _GEN_2396;
        end else begin
          tag_87 <= _GEN_4723;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_88 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_88 <= _GEN_2397;
        end else begin
          tag_88 <= _GEN_4724;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_89 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_89 <= _GEN_2398;
        end else begin
          tag_89 <= _GEN_4725;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_90 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_90 <= _GEN_2399;
        end else begin
          tag_90 <= _GEN_4726;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_91 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_91 <= _GEN_2400;
        end else begin
          tag_91 <= _GEN_4727;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_92 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_92 <= _GEN_2401;
        end else begin
          tag_92 <= _GEN_4728;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_93 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_93 <= _GEN_2402;
        end else begin
          tag_93 <= _GEN_4729;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_94 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_94 <= _GEN_2403;
        end else begin
          tag_94 <= _GEN_4730;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_95 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_95 <= _GEN_2404;
        end else begin
          tag_95 <= _GEN_4731;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_96 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_96 <= _GEN_2405;
        end else begin
          tag_96 <= _GEN_4732;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_97 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_97 <= _GEN_2406;
        end else begin
          tag_97 <= _GEN_4733;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_98 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_98 <= _GEN_2407;
        end else begin
          tag_98 <= _GEN_4734;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_99 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_99 <= _GEN_2408;
        end else begin
          tag_99 <= _GEN_4735;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_100 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_100 <= _GEN_2409;
        end else begin
          tag_100 <= _GEN_4736;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_101 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_101 <= _GEN_2410;
        end else begin
          tag_101 <= _GEN_4737;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_102 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_102 <= _GEN_2411;
        end else begin
          tag_102 <= _GEN_4738;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_103 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_103 <= _GEN_2412;
        end else begin
          tag_103 <= _GEN_4739;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_104 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_104 <= _GEN_2413;
        end else begin
          tag_104 <= _GEN_4740;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_105 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_105 <= _GEN_2414;
        end else begin
          tag_105 <= _GEN_4741;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_106 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_106 <= _GEN_2415;
        end else begin
          tag_106 <= _GEN_4742;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_107 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_107 <= _GEN_2416;
        end else begin
          tag_107 <= _GEN_4743;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_108 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_108 <= _GEN_2417;
        end else begin
          tag_108 <= _GEN_4744;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_109 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_109 <= _GEN_2418;
        end else begin
          tag_109 <= _GEN_4745;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_110 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_110 <= _GEN_2419;
        end else begin
          tag_110 <= _GEN_4746;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_111 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_111 <= _GEN_2420;
        end else begin
          tag_111 <= _GEN_4747;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_112 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_112 <= _GEN_2421;
        end else begin
          tag_112 <= _GEN_4748;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_113 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_113 <= _GEN_2422;
        end else begin
          tag_113 <= _GEN_4749;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_114 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_114 <= _GEN_2423;
        end else begin
          tag_114 <= _GEN_4750;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_115 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_115 <= _GEN_2424;
        end else begin
          tag_115 <= _GEN_4751;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_116 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_116 <= _GEN_2425;
        end else begin
          tag_116 <= _GEN_4752;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_117 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_117 <= _GEN_2426;
        end else begin
          tag_117 <= _GEN_4753;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_118 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_118 <= _GEN_2427;
        end else begin
          tag_118 <= _GEN_4754;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_119 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_119 <= _GEN_2428;
        end else begin
          tag_119 <= _GEN_4755;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_120 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_120 <= _GEN_2429;
        end else begin
          tag_120 <= _GEN_4756;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_121 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_121 <= _GEN_2430;
        end else begin
          tag_121 <= _GEN_4757;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_122 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_122 <= _GEN_2431;
        end else begin
          tag_122 <= _GEN_4758;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_123 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_123 <= _GEN_2432;
        end else begin
          tag_123 <= _GEN_4759;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_124 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_124 <= _GEN_2433;
        end else begin
          tag_124 <= _GEN_4760;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_125 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_125 <= _GEN_2434;
        end else begin
          tag_125 <= _GEN_4761;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_126 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_126 <= _GEN_2435;
        end else begin
          tag_126 <= _GEN_4762;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_127 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_127 <= _GEN_2436;
        end else begin
          tag_127 <= _GEN_4763;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_128 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_128 <= _GEN_2437;
        end else begin
          tag_128 <= _GEN_4764;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_129 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_129 <= _GEN_2438;
        end else begin
          tag_129 <= _GEN_4765;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_130 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_130 <= _GEN_2439;
        end else begin
          tag_130 <= _GEN_4766;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_131 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_131 <= _GEN_2440;
        end else begin
          tag_131 <= _GEN_4767;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_132 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_132 <= _GEN_2441;
        end else begin
          tag_132 <= _GEN_4768;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_133 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_133 <= _GEN_2442;
        end else begin
          tag_133 <= _GEN_4769;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_134 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_134 <= _GEN_2443;
        end else begin
          tag_134 <= _GEN_4770;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_135 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_135 <= _GEN_2444;
        end else begin
          tag_135 <= _GEN_4771;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_136 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_136 <= _GEN_2445;
        end else begin
          tag_136 <= _GEN_4772;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_137 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_137 <= _GEN_2446;
        end else begin
          tag_137 <= _GEN_4773;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_138 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_138 <= _GEN_2447;
        end else begin
          tag_138 <= _GEN_4774;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_139 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_139 <= _GEN_2448;
        end else begin
          tag_139 <= _GEN_4775;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_140 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_140 <= _GEN_2449;
        end else begin
          tag_140 <= _GEN_4776;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_141 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_141 <= _GEN_2450;
        end else begin
          tag_141 <= _GEN_4777;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_142 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_142 <= _GEN_2451;
        end else begin
          tag_142 <= _GEN_4778;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_143 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_143 <= _GEN_2452;
        end else begin
          tag_143 <= _GEN_4779;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_144 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_144 <= _GEN_2453;
        end else begin
          tag_144 <= _GEN_4780;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_145 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_145 <= _GEN_2454;
        end else begin
          tag_145 <= _GEN_4781;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_146 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_146 <= _GEN_2455;
        end else begin
          tag_146 <= _GEN_4782;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_147 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_147 <= _GEN_2456;
        end else begin
          tag_147 <= _GEN_4783;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_148 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_148 <= _GEN_2457;
        end else begin
          tag_148 <= _GEN_4784;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_149 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_149 <= _GEN_2458;
        end else begin
          tag_149 <= _GEN_4785;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_150 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_150 <= _GEN_2459;
        end else begin
          tag_150 <= _GEN_4786;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_151 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_151 <= _GEN_2460;
        end else begin
          tag_151 <= _GEN_4787;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_152 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_152 <= _GEN_2461;
        end else begin
          tag_152 <= _GEN_4788;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_153 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_153 <= _GEN_2462;
        end else begin
          tag_153 <= _GEN_4789;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_154 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_154 <= _GEN_2463;
        end else begin
          tag_154 <= _GEN_4790;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_155 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_155 <= _GEN_2464;
        end else begin
          tag_155 <= _GEN_4791;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_156 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_156 <= _GEN_2465;
        end else begin
          tag_156 <= _GEN_4792;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_157 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_157 <= _GEN_2466;
        end else begin
          tag_157 <= _GEN_4793;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_158 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_158 <= _GEN_2467;
        end else begin
          tag_158 <= _GEN_4794;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_159 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_159 <= _GEN_2468;
        end else begin
          tag_159 <= _GEN_4795;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_160 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_160 <= _GEN_2469;
        end else begin
          tag_160 <= _GEN_4796;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_161 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_161 <= _GEN_2470;
        end else begin
          tag_161 <= _GEN_4797;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_162 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_162 <= _GEN_2471;
        end else begin
          tag_162 <= _GEN_4798;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_163 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_163 <= _GEN_2472;
        end else begin
          tag_163 <= _GEN_4799;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_164 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_164 <= _GEN_2473;
        end else begin
          tag_164 <= _GEN_4800;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_165 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_165 <= _GEN_2474;
        end else begin
          tag_165 <= _GEN_4801;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_166 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_166 <= _GEN_2475;
        end else begin
          tag_166 <= _GEN_4802;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_167 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_167 <= _GEN_2476;
        end else begin
          tag_167 <= _GEN_4803;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_168 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_168 <= _GEN_2477;
        end else begin
          tag_168 <= _GEN_4804;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_169 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_169 <= _GEN_2478;
        end else begin
          tag_169 <= _GEN_4805;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_170 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_170 <= _GEN_2479;
        end else begin
          tag_170 <= _GEN_4806;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_171 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_171 <= _GEN_2480;
        end else begin
          tag_171 <= _GEN_4807;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_172 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_172 <= _GEN_2481;
        end else begin
          tag_172 <= _GEN_4808;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_173 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_173 <= _GEN_2482;
        end else begin
          tag_173 <= _GEN_4809;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_174 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_174 <= _GEN_2483;
        end else begin
          tag_174 <= _GEN_4810;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_175 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_175 <= _GEN_2484;
        end else begin
          tag_175 <= _GEN_4811;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_176 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_176 <= _GEN_2485;
        end else begin
          tag_176 <= _GEN_4812;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_177 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_177 <= _GEN_2486;
        end else begin
          tag_177 <= _GEN_4813;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_178 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_178 <= _GEN_2487;
        end else begin
          tag_178 <= _GEN_4814;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_179 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_179 <= _GEN_2488;
        end else begin
          tag_179 <= _GEN_4815;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_180 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_180 <= _GEN_2489;
        end else begin
          tag_180 <= _GEN_4816;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_181 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_181 <= _GEN_2490;
        end else begin
          tag_181 <= _GEN_4817;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_182 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_182 <= _GEN_2491;
        end else begin
          tag_182 <= _GEN_4818;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_183 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_183 <= _GEN_2492;
        end else begin
          tag_183 <= _GEN_4819;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_184 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_184 <= _GEN_2493;
        end else begin
          tag_184 <= _GEN_4820;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_185 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_185 <= _GEN_2494;
        end else begin
          tag_185 <= _GEN_4821;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_186 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_186 <= _GEN_2495;
        end else begin
          tag_186 <= _GEN_4822;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_187 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_187 <= _GEN_2496;
        end else begin
          tag_187 <= _GEN_4823;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_188 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_188 <= _GEN_2497;
        end else begin
          tag_188 <= _GEN_4824;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_189 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_189 <= _GEN_2498;
        end else begin
          tag_189 <= _GEN_4825;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_190 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_190 <= _GEN_2499;
        end else begin
          tag_190 <= _GEN_4826;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_191 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_191 <= _GEN_2500;
        end else begin
          tag_191 <= _GEN_4827;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_192 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_192 <= _GEN_2501;
        end else begin
          tag_192 <= _GEN_4828;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_193 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_193 <= _GEN_2502;
        end else begin
          tag_193 <= _GEN_4829;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_194 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_194 <= _GEN_2503;
        end else begin
          tag_194 <= _GEN_4830;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_195 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_195 <= _GEN_2504;
        end else begin
          tag_195 <= _GEN_4831;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_196 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_196 <= _GEN_2505;
        end else begin
          tag_196 <= _GEN_4832;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_197 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_197 <= _GEN_2506;
        end else begin
          tag_197 <= _GEN_4833;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_198 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_198 <= _GEN_2507;
        end else begin
          tag_198 <= _GEN_4834;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_199 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_199 <= _GEN_2508;
        end else begin
          tag_199 <= _GEN_4835;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_200 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_200 <= _GEN_2509;
        end else begin
          tag_200 <= _GEN_4836;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_201 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_201 <= _GEN_2510;
        end else begin
          tag_201 <= _GEN_4837;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_202 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_202 <= _GEN_2511;
        end else begin
          tag_202 <= _GEN_4838;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_203 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_203 <= _GEN_2512;
        end else begin
          tag_203 <= _GEN_4839;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_204 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_204 <= _GEN_2513;
        end else begin
          tag_204 <= _GEN_4840;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_205 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_205 <= _GEN_2514;
        end else begin
          tag_205 <= _GEN_4841;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_206 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_206 <= _GEN_2515;
        end else begin
          tag_206 <= _GEN_4842;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_207 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_207 <= _GEN_2516;
        end else begin
          tag_207 <= _GEN_4843;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_208 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_208 <= _GEN_2517;
        end else begin
          tag_208 <= _GEN_4844;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_209 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_209 <= _GEN_2518;
        end else begin
          tag_209 <= _GEN_4845;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_210 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_210 <= _GEN_2519;
        end else begin
          tag_210 <= _GEN_4846;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_211 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_211 <= _GEN_2520;
        end else begin
          tag_211 <= _GEN_4847;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_212 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_212 <= _GEN_2521;
        end else begin
          tag_212 <= _GEN_4848;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_213 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_213 <= _GEN_2522;
        end else begin
          tag_213 <= _GEN_4849;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_214 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_214 <= _GEN_2523;
        end else begin
          tag_214 <= _GEN_4850;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_215 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_215 <= _GEN_2524;
        end else begin
          tag_215 <= _GEN_4851;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_216 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_216 <= _GEN_2525;
        end else begin
          tag_216 <= _GEN_4852;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_217 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_217 <= _GEN_2526;
        end else begin
          tag_217 <= _GEN_4853;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_218 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_218 <= _GEN_2527;
        end else begin
          tag_218 <= _GEN_4854;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_219 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_219 <= _GEN_2528;
        end else begin
          tag_219 <= _GEN_4855;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_220 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_220 <= _GEN_2529;
        end else begin
          tag_220 <= _GEN_4856;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_221 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_221 <= _GEN_2530;
        end else begin
          tag_221 <= _GEN_4857;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_222 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_222 <= _GEN_2531;
        end else begin
          tag_222 <= _GEN_4858;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_223 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_223 <= _GEN_2532;
        end else begin
          tag_223 <= _GEN_4859;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_224 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_224 <= _GEN_2533;
        end else begin
          tag_224 <= _GEN_4860;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_225 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_225 <= _GEN_2534;
        end else begin
          tag_225 <= _GEN_4861;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_226 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_226 <= _GEN_2535;
        end else begin
          tag_226 <= _GEN_4862;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_227 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_227 <= _GEN_2536;
        end else begin
          tag_227 <= _GEN_4863;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_228 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_228 <= _GEN_2537;
        end else begin
          tag_228 <= _GEN_4864;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_229 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_229 <= _GEN_2538;
        end else begin
          tag_229 <= _GEN_4865;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_230 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_230 <= _GEN_2539;
        end else begin
          tag_230 <= _GEN_4866;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_231 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_231 <= _GEN_2540;
        end else begin
          tag_231 <= _GEN_4867;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_232 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_232 <= _GEN_2541;
        end else begin
          tag_232 <= _GEN_4868;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_233 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_233 <= _GEN_2542;
        end else begin
          tag_233 <= _GEN_4869;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_234 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_234 <= _GEN_2543;
        end else begin
          tag_234 <= _GEN_4870;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_235 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_235 <= _GEN_2544;
        end else begin
          tag_235 <= _GEN_4871;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_236 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_236 <= _GEN_2545;
        end else begin
          tag_236 <= _GEN_4872;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_237 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_237 <= _GEN_2546;
        end else begin
          tag_237 <= _GEN_4873;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_238 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_238 <= _GEN_2547;
        end else begin
          tag_238 <= _GEN_4874;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_239 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_239 <= _GEN_2548;
        end else begin
          tag_239 <= _GEN_4875;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_240 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_240 <= _GEN_2549;
        end else begin
          tag_240 <= _GEN_4876;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_241 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_241 <= _GEN_2550;
        end else begin
          tag_241 <= _GEN_4877;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_242 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_242 <= _GEN_2551;
        end else begin
          tag_242 <= _GEN_4878;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_243 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_243 <= _GEN_2552;
        end else begin
          tag_243 <= _GEN_4879;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_244 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_244 <= _GEN_2553;
        end else begin
          tag_244 <= _GEN_4880;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_245 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_245 <= _GEN_2554;
        end else begin
          tag_245 <= _GEN_4881;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_246 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_246 <= _GEN_2555;
        end else begin
          tag_246 <= _GEN_4882;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_247 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_247 <= _GEN_2556;
        end else begin
          tag_247 <= _GEN_4883;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_248 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_248 <= _GEN_2557;
        end else begin
          tag_248 <= _GEN_4884;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_249 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_249 <= _GEN_2558;
        end else begin
          tag_249 <= _GEN_4885;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_250 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_250 <= _GEN_2559;
        end else begin
          tag_250 <= _GEN_4886;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_251 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_251 <= _GEN_2560;
        end else begin
          tag_251 <= _GEN_4887;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_252 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_252 <= _GEN_2561;
        end else begin
          tag_252 <= _GEN_4888;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_253 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_253 <= _GEN_2562;
        end else begin
          tag_253 <= _GEN_4889;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_254 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_254 <= _GEN_2563;
        end else begin
          tag_254 <= _GEN_4890;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      tag_255 <= 20'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          tag_255 <= _GEN_2564;
        end else begin
          tag_255 <= _GEN_4891;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_0 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_0 <= _GEN_2053;
        end else begin
          valid_0 <= _GEN_4380;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_1 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_1 <= _GEN_2054;
        end else begin
          valid_1 <= _GEN_4381;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_2 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_2 <= _GEN_2055;
        end else begin
          valid_2 <= _GEN_4382;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_3 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_3 <= _GEN_2056;
        end else begin
          valid_3 <= _GEN_4383;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_4 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_4 <= _GEN_2057;
        end else begin
          valid_4 <= _GEN_4384;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_5 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_5 <= _GEN_2058;
        end else begin
          valid_5 <= _GEN_4385;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_6 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_6 <= _GEN_2059;
        end else begin
          valid_6 <= _GEN_4386;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_7 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_7 <= _GEN_2060;
        end else begin
          valid_7 <= _GEN_4387;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_8 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_8 <= _GEN_2061;
        end else begin
          valid_8 <= _GEN_4388;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_9 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_9 <= _GEN_2062;
        end else begin
          valid_9 <= _GEN_4389;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_10 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_10 <= _GEN_2063;
        end else begin
          valid_10 <= _GEN_4390;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_11 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_11 <= _GEN_2064;
        end else begin
          valid_11 <= _GEN_4391;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_12 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_12 <= _GEN_2065;
        end else begin
          valid_12 <= _GEN_4392;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_13 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_13 <= _GEN_2066;
        end else begin
          valid_13 <= _GEN_4393;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_14 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_14 <= _GEN_2067;
        end else begin
          valid_14 <= _GEN_4394;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_15 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_15 <= _GEN_2068;
        end else begin
          valid_15 <= _GEN_4395;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_16 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_16 <= _GEN_2069;
        end else begin
          valid_16 <= _GEN_4396;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_17 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_17 <= _GEN_2070;
        end else begin
          valid_17 <= _GEN_4397;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_18 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_18 <= _GEN_2071;
        end else begin
          valid_18 <= _GEN_4398;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_19 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_19 <= _GEN_2072;
        end else begin
          valid_19 <= _GEN_4399;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_20 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_20 <= _GEN_2073;
        end else begin
          valid_20 <= _GEN_4400;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_21 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_21 <= _GEN_2074;
        end else begin
          valid_21 <= _GEN_4401;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_22 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_22 <= _GEN_2075;
        end else begin
          valid_22 <= _GEN_4402;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_23 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_23 <= _GEN_2076;
        end else begin
          valid_23 <= _GEN_4403;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_24 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_24 <= _GEN_2077;
        end else begin
          valid_24 <= _GEN_4404;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_25 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_25 <= _GEN_2078;
        end else begin
          valid_25 <= _GEN_4405;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_26 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_26 <= _GEN_2079;
        end else begin
          valid_26 <= _GEN_4406;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_27 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_27 <= _GEN_2080;
        end else begin
          valid_27 <= _GEN_4407;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_28 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_28 <= _GEN_2081;
        end else begin
          valid_28 <= _GEN_4408;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_29 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_29 <= _GEN_2082;
        end else begin
          valid_29 <= _GEN_4409;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_30 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_30 <= _GEN_2083;
        end else begin
          valid_30 <= _GEN_4410;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_31 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_31 <= _GEN_2084;
        end else begin
          valid_31 <= _GEN_4411;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_32 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_32 <= _GEN_2085;
        end else begin
          valid_32 <= _GEN_4412;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_33 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_33 <= _GEN_2086;
        end else begin
          valid_33 <= _GEN_4413;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_34 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_34 <= _GEN_2087;
        end else begin
          valid_34 <= _GEN_4414;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_35 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_35 <= _GEN_2088;
        end else begin
          valid_35 <= _GEN_4415;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_36 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_36 <= _GEN_2089;
        end else begin
          valid_36 <= _GEN_4416;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_37 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_37 <= _GEN_2090;
        end else begin
          valid_37 <= _GEN_4417;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_38 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_38 <= _GEN_2091;
        end else begin
          valid_38 <= _GEN_4418;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_39 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_39 <= _GEN_2092;
        end else begin
          valid_39 <= _GEN_4419;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_40 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_40 <= _GEN_2093;
        end else begin
          valid_40 <= _GEN_4420;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_41 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_41 <= _GEN_2094;
        end else begin
          valid_41 <= _GEN_4421;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_42 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_42 <= _GEN_2095;
        end else begin
          valid_42 <= _GEN_4422;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_43 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_43 <= _GEN_2096;
        end else begin
          valid_43 <= _GEN_4423;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_44 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_44 <= _GEN_2097;
        end else begin
          valid_44 <= _GEN_4424;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_45 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_45 <= _GEN_2098;
        end else begin
          valid_45 <= _GEN_4425;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_46 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_46 <= _GEN_2099;
        end else begin
          valid_46 <= _GEN_4426;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_47 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_47 <= _GEN_2100;
        end else begin
          valid_47 <= _GEN_4427;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_48 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_48 <= _GEN_2101;
        end else begin
          valid_48 <= _GEN_4428;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_49 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_49 <= _GEN_2102;
        end else begin
          valid_49 <= _GEN_4429;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_50 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_50 <= _GEN_2103;
        end else begin
          valid_50 <= _GEN_4430;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_51 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_51 <= _GEN_2104;
        end else begin
          valid_51 <= _GEN_4431;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_52 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_52 <= _GEN_2105;
        end else begin
          valid_52 <= _GEN_4432;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_53 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_53 <= _GEN_2106;
        end else begin
          valid_53 <= _GEN_4433;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_54 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_54 <= _GEN_2107;
        end else begin
          valid_54 <= _GEN_4434;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_55 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_55 <= _GEN_2108;
        end else begin
          valid_55 <= _GEN_4435;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_56 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_56 <= _GEN_2109;
        end else begin
          valid_56 <= _GEN_4436;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_57 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_57 <= _GEN_2110;
        end else begin
          valid_57 <= _GEN_4437;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_58 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_58 <= _GEN_2111;
        end else begin
          valid_58 <= _GEN_4438;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_59 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_59 <= _GEN_2112;
        end else begin
          valid_59 <= _GEN_4439;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_60 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_60 <= _GEN_2113;
        end else begin
          valid_60 <= _GEN_4440;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_61 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_61 <= _GEN_2114;
        end else begin
          valid_61 <= _GEN_4441;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_62 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_62 <= _GEN_2115;
        end else begin
          valid_62 <= _GEN_4442;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_63 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_63 <= _GEN_2116;
        end else begin
          valid_63 <= _GEN_4443;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_64 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_64 <= _GEN_2117;
        end else begin
          valid_64 <= _GEN_4444;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_65 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_65 <= _GEN_2118;
        end else begin
          valid_65 <= _GEN_4445;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_66 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_66 <= _GEN_2119;
        end else begin
          valid_66 <= _GEN_4446;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_67 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_67 <= _GEN_2120;
        end else begin
          valid_67 <= _GEN_4447;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_68 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_68 <= _GEN_2121;
        end else begin
          valid_68 <= _GEN_4448;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_69 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_69 <= _GEN_2122;
        end else begin
          valid_69 <= _GEN_4449;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_70 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_70 <= _GEN_2123;
        end else begin
          valid_70 <= _GEN_4450;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_71 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_71 <= _GEN_2124;
        end else begin
          valid_71 <= _GEN_4451;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_72 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_72 <= _GEN_2125;
        end else begin
          valid_72 <= _GEN_4452;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_73 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_73 <= _GEN_2126;
        end else begin
          valid_73 <= _GEN_4453;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_74 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_74 <= _GEN_2127;
        end else begin
          valid_74 <= _GEN_4454;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_75 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_75 <= _GEN_2128;
        end else begin
          valid_75 <= _GEN_4455;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_76 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_76 <= _GEN_2129;
        end else begin
          valid_76 <= _GEN_4456;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_77 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_77 <= _GEN_2130;
        end else begin
          valid_77 <= _GEN_4457;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_78 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_78 <= _GEN_2131;
        end else begin
          valid_78 <= _GEN_4458;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_79 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_79 <= _GEN_2132;
        end else begin
          valid_79 <= _GEN_4459;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_80 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_80 <= _GEN_2133;
        end else begin
          valid_80 <= _GEN_4460;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_81 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_81 <= _GEN_2134;
        end else begin
          valid_81 <= _GEN_4461;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_82 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_82 <= _GEN_2135;
        end else begin
          valid_82 <= _GEN_4462;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_83 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_83 <= _GEN_2136;
        end else begin
          valid_83 <= _GEN_4463;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_84 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_84 <= _GEN_2137;
        end else begin
          valid_84 <= _GEN_4464;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_85 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_85 <= _GEN_2138;
        end else begin
          valid_85 <= _GEN_4465;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_86 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_86 <= _GEN_2139;
        end else begin
          valid_86 <= _GEN_4466;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_87 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_87 <= _GEN_2140;
        end else begin
          valid_87 <= _GEN_4467;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_88 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_88 <= _GEN_2141;
        end else begin
          valid_88 <= _GEN_4468;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_89 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_89 <= _GEN_2142;
        end else begin
          valid_89 <= _GEN_4469;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_90 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_90 <= _GEN_2143;
        end else begin
          valid_90 <= _GEN_4470;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_91 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_91 <= _GEN_2144;
        end else begin
          valid_91 <= _GEN_4471;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_92 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_92 <= _GEN_2145;
        end else begin
          valid_92 <= _GEN_4472;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_93 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_93 <= _GEN_2146;
        end else begin
          valid_93 <= _GEN_4473;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_94 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_94 <= _GEN_2147;
        end else begin
          valid_94 <= _GEN_4474;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_95 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_95 <= _GEN_2148;
        end else begin
          valid_95 <= _GEN_4475;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_96 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_96 <= _GEN_2149;
        end else begin
          valid_96 <= _GEN_4476;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_97 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_97 <= _GEN_2150;
        end else begin
          valid_97 <= _GEN_4477;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_98 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_98 <= _GEN_2151;
        end else begin
          valid_98 <= _GEN_4478;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_99 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_99 <= _GEN_2152;
        end else begin
          valid_99 <= _GEN_4479;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_100 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_100 <= _GEN_2153;
        end else begin
          valid_100 <= _GEN_4480;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_101 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_101 <= _GEN_2154;
        end else begin
          valid_101 <= _GEN_4481;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_102 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_102 <= _GEN_2155;
        end else begin
          valid_102 <= _GEN_4482;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_103 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_103 <= _GEN_2156;
        end else begin
          valid_103 <= _GEN_4483;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_104 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_104 <= _GEN_2157;
        end else begin
          valid_104 <= _GEN_4484;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_105 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_105 <= _GEN_2158;
        end else begin
          valid_105 <= _GEN_4485;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_106 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_106 <= _GEN_2159;
        end else begin
          valid_106 <= _GEN_4486;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_107 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_107 <= _GEN_2160;
        end else begin
          valid_107 <= _GEN_4487;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_108 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_108 <= _GEN_2161;
        end else begin
          valid_108 <= _GEN_4488;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_109 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_109 <= _GEN_2162;
        end else begin
          valid_109 <= _GEN_4489;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_110 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_110 <= _GEN_2163;
        end else begin
          valid_110 <= _GEN_4490;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_111 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_111 <= _GEN_2164;
        end else begin
          valid_111 <= _GEN_4491;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_112 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_112 <= _GEN_2165;
        end else begin
          valid_112 <= _GEN_4492;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_113 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_113 <= _GEN_2166;
        end else begin
          valid_113 <= _GEN_4493;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_114 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_114 <= _GEN_2167;
        end else begin
          valid_114 <= _GEN_4494;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_115 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_115 <= _GEN_2168;
        end else begin
          valid_115 <= _GEN_4495;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_116 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_116 <= _GEN_2169;
        end else begin
          valid_116 <= _GEN_4496;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_117 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_117 <= _GEN_2170;
        end else begin
          valid_117 <= _GEN_4497;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_118 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_118 <= _GEN_2171;
        end else begin
          valid_118 <= _GEN_4498;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_119 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_119 <= _GEN_2172;
        end else begin
          valid_119 <= _GEN_4499;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_120 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_120 <= _GEN_2173;
        end else begin
          valid_120 <= _GEN_4500;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_121 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_121 <= _GEN_2174;
        end else begin
          valid_121 <= _GEN_4501;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_122 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_122 <= _GEN_2175;
        end else begin
          valid_122 <= _GEN_4502;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_123 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_123 <= _GEN_2176;
        end else begin
          valid_123 <= _GEN_4503;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_124 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_124 <= _GEN_2177;
        end else begin
          valid_124 <= _GEN_4504;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_125 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_125 <= _GEN_2178;
        end else begin
          valid_125 <= _GEN_4505;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_126 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_126 <= _GEN_2179;
        end else begin
          valid_126 <= _GEN_4506;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_127 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_127 <= _GEN_2180;
        end else begin
          valid_127 <= _GEN_4507;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_128 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_128 <= _GEN_2181;
        end else begin
          valid_128 <= _GEN_4508;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_129 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_129 <= _GEN_2182;
        end else begin
          valid_129 <= _GEN_4509;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_130 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_130 <= _GEN_2183;
        end else begin
          valid_130 <= _GEN_4510;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_131 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_131 <= _GEN_2184;
        end else begin
          valid_131 <= _GEN_4511;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_132 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_132 <= _GEN_2185;
        end else begin
          valid_132 <= _GEN_4512;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_133 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_133 <= _GEN_2186;
        end else begin
          valid_133 <= _GEN_4513;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_134 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_134 <= _GEN_2187;
        end else begin
          valid_134 <= _GEN_4514;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_135 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_135 <= _GEN_2188;
        end else begin
          valid_135 <= _GEN_4515;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_136 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_136 <= _GEN_2189;
        end else begin
          valid_136 <= _GEN_4516;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_137 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_137 <= _GEN_2190;
        end else begin
          valid_137 <= _GEN_4517;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_138 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_138 <= _GEN_2191;
        end else begin
          valid_138 <= _GEN_4518;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_139 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_139 <= _GEN_2192;
        end else begin
          valid_139 <= _GEN_4519;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_140 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_140 <= _GEN_2193;
        end else begin
          valid_140 <= _GEN_4520;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_141 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_141 <= _GEN_2194;
        end else begin
          valid_141 <= _GEN_4521;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_142 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_142 <= _GEN_2195;
        end else begin
          valid_142 <= _GEN_4522;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_143 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_143 <= _GEN_2196;
        end else begin
          valid_143 <= _GEN_4523;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_144 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_144 <= _GEN_2197;
        end else begin
          valid_144 <= _GEN_4524;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_145 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_145 <= _GEN_2198;
        end else begin
          valid_145 <= _GEN_4525;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_146 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_146 <= _GEN_2199;
        end else begin
          valid_146 <= _GEN_4526;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_147 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_147 <= _GEN_2200;
        end else begin
          valid_147 <= _GEN_4527;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_148 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_148 <= _GEN_2201;
        end else begin
          valid_148 <= _GEN_4528;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_149 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_149 <= _GEN_2202;
        end else begin
          valid_149 <= _GEN_4529;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_150 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_150 <= _GEN_2203;
        end else begin
          valid_150 <= _GEN_4530;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_151 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_151 <= _GEN_2204;
        end else begin
          valid_151 <= _GEN_4531;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_152 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_152 <= _GEN_2205;
        end else begin
          valid_152 <= _GEN_4532;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_153 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_153 <= _GEN_2206;
        end else begin
          valid_153 <= _GEN_4533;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_154 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_154 <= _GEN_2207;
        end else begin
          valid_154 <= _GEN_4534;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_155 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_155 <= _GEN_2208;
        end else begin
          valid_155 <= _GEN_4535;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_156 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_156 <= _GEN_2209;
        end else begin
          valid_156 <= _GEN_4536;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_157 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_157 <= _GEN_2210;
        end else begin
          valid_157 <= _GEN_4537;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_158 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_158 <= _GEN_2211;
        end else begin
          valid_158 <= _GEN_4538;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_159 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_159 <= _GEN_2212;
        end else begin
          valid_159 <= _GEN_4539;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_160 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_160 <= _GEN_2213;
        end else begin
          valid_160 <= _GEN_4540;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_161 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_161 <= _GEN_2214;
        end else begin
          valid_161 <= _GEN_4541;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_162 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_162 <= _GEN_2215;
        end else begin
          valid_162 <= _GEN_4542;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_163 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_163 <= _GEN_2216;
        end else begin
          valid_163 <= _GEN_4543;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_164 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_164 <= _GEN_2217;
        end else begin
          valid_164 <= _GEN_4544;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_165 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_165 <= _GEN_2218;
        end else begin
          valid_165 <= _GEN_4545;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_166 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_166 <= _GEN_2219;
        end else begin
          valid_166 <= _GEN_4546;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_167 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_167 <= _GEN_2220;
        end else begin
          valid_167 <= _GEN_4547;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_168 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_168 <= _GEN_2221;
        end else begin
          valid_168 <= _GEN_4548;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_169 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_169 <= _GEN_2222;
        end else begin
          valid_169 <= _GEN_4549;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_170 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_170 <= _GEN_2223;
        end else begin
          valid_170 <= _GEN_4550;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_171 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_171 <= _GEN_2224;
        end else begin
          valid_171 <= _GEN_4551;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_172 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_172 <= _GEN_2225;
        end else begin
          valid_172 <= _GEN_4552;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_173 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_173 <= _GEN_2226;
        end else begin
          valid_173 <= _GEN_4553;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_174 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_174 <= _GEN_2227;
        end else begin
          valid_174 <= _GEN_4554;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_175 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_175 <= _GEN_2228;
        end else begin
          valid_175 <= _GEN_4555;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_176 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_176 <= _GEN_2229;
        end else begin
          valid_176 <= _GEN_4556;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_177 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_177 <= _GEN_2230;
        end else begin
          valid_177 <= _GEN_4557;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_178 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_178 <= _GEN_2231;
        end else begin
          valid_178 <= _GEN_4558;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_179 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_179 <= _GEN_2232;
        end else begin
          valid_179 <= _GEN_4559;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_180 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_180 <= _GEN_2233;
        end else begin
          valid_180 <= _GEN_4560;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_181 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_181 <= _GEN_2234;
        end else begin
          valid_181 <= _GEN_4561;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_182 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_182 <= _GEN_2235;
        end else begin
          valid_182 <= _GEN_4562;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_183 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_183 <= _GEN_2236;
        end else begin
          valid_183 <= _GEN_4563;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_184 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_184 <= _GEN_2237;
        end else begin
          valid_184 <= _GEN_4564;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_185 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_185 <= _GEN_2238;
        end else begin
          valid_185 <= _GEN_4565;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_186 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_186 <= _GEN_2239;
        end else begin
          valid_186 <= _GEN_4566;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_187 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_187 <= _GEN_2240;
        end else begin
          valid_187 <= _GEN_4567;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_188 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_188 <= _GEN_2241;
        end else begin
          valid_188 <= _GEN_4568;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_189 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_189 <= _GEN_2242;
        end else begin
          valid_189 <= _GEN_4569;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_190 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_190 <= _GEN_2243;
        end else begin
          valid_190 <= _GEN_4570;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_191 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_191 <= _GEN_2244;
        end else begin
          valid_191 <= _GEN_4571;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_192 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_192 <= _GEN_2245;
        end else begin
          valid_192 <= _GEN_4572;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_193 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_193 <= _GEN_2246;
        end else begin
          valid_193 <= _GEN_4573;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_194 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_194 <= _GEN_2247;
        end else begin
          valid_194 <= _GEN_4574;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_195 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_195 <= _GEN_2248;
        end else begin
          valid_195 <= _GEN_4575;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_196 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_196 <= _GEN_2249;
        end else begin
          valid_196 <= _GEN_4576;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_197 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_197 <= _GEN_2250;
        end else begin
          valid_197 <= _GEN_4577;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_198 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_198 <= _GEN_2251;
        end else begin
          valid_198 <= _GEN_4578;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_199 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_199 <= _GEN_2252;
        end else begin
          valid_199 <= _GEN_4579;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_200 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_200 <= _GEN_2253;
        end else begin
          valid_200 <= _GEN_4580;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_201 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_201 <= _GEN_2254;
        end else begin
          valid_201 <= _GEN_4581;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_202 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_202 <= _GEN_2255;
        end else begin
          valid_202 <= _GEN_4582;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_203 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_203 <= _GEN_2256;
        end else begin
          valid_203 <= _GEN_4583;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_204 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_204 <= _GEN_2257;
        end else begin
          valid_204 <= _GEN_4584;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_205 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_205 <= _GEN_2258;
        end else begin
          valid_205 <= _GEN_4585;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_206 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_206 <= _GEN_2259;
        end else begin
          valid_206 <= _GEN_4586;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_207 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_207 <= _GEN_2260;
        end else begin
          valid_207 <= _GEN_4587;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_208 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_208 <= _GEN_2261;
        end else begin
          valid_208 <= _GEN_4588;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_209 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_209 <= _GEN_2262;
        end else begin
          valid_209 <= _GEN_4589;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_210 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_210 <= _GEN_2263;
        end else begin
          valid_210 <= _GEN_4590;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_211 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_211 <= _GEN_2264;
        end else begin
          valid_211 <= _GEN_4591;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_212 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_212 <= _GEN_2265;
        end else begin
          valid_212 <= _GEN_4592;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_213 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_213 <= _GEN_2266;
        end else begin
          valid_213 <= _GEN_4593;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_214 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_214 <= _GEN_2267;
        end else begin
          valid_214 <= _GEN_4594;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_215 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_215 <= _GEN_2268;
        end else begin
          valid_215 <= _GEN_4595;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_216 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_216 <= _GEN_2269;
        end else begin
          valid_216 <= _GEN_4596;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_217 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_217 <= _GEN_2270;
        end else begin
          valid_217 <= _GEN_4597;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_218 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_218 <= _GEN_2271;
        end else begin
          valid_218 <= _GEN_4598;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_219 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_219 <= _GEN_2272;
        end else begin
          valid_219 <= _GEN_4599;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_220 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_220 <= _GEN_2273;
        end else begin
          valid_220 <= _GEN_4600;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_221 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_221 <= _GEN_2274;
        end else begin
          valid_221 <= _GEN_4601;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_222 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_222 <= _GEN_2275;
        end else begin
          valid_222 <= _GEN_4602;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_223 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_223 <= _GEN_2276;
        end else begin
          valid_223 <= _GEN_4603;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_224 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_224 <= _GEN_2277;
        end else begin
          valid_224 <= _GEN_4604;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_225 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_225 <= _GEN_2278;
        end else begin
          valid_225 <= _GEN_4605;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_226 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_226 <= _GEN_2279;
        end else begin
          valid_226 <= _GEN_4606;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_227 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_227 <= _GEN_2280;
        end else begin
          valid_227 <= _GEN_4607;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_228 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_228 <= _GEN_2281;
        end else begin
          valid_228 <= _GEN_4608;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_229 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_229 <= _GEN_2282;
        end else begin
          valid_229 <= _GEN_4609;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_230 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_230 <= _GEN_2283;
        end else begin
          valid_230 <= _GEN_4610;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_231 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_231 <= _GEN_2284;
        end else begin
          valid_231 <= _GEN_4611;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_232 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_232 <= _GEN_2285;
        end else begin
          valid_232 <= _GEN_4612;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_233 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_233 <= _GEN_2286;
        end else begin
          valid_233 <= _GEN_4613;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_234 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_234 <= _GEN_2287;
        end else begin
          valid_234 <= _GEN_4614;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_235 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_235 <= _GEN_2288;
        end else begin
          valid_235 <= _GEN_4615;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_236 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_236 <= _GEN_2289;
        end else begin
          valid_236 <= _GEN_4616;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_237 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_237 <= _GEN_2290;
        end else begin
          valid_237 <= _GEN_4617;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_238 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_238 <= _GEN_2291;
        end else begin
          valid_238 <= _GEN_4618;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_239 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_239 <= _GEN_2292;
        end else begin
          valid_239 <= _GEN_4619;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_240 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_240 <= _GEN_2293;
        end else begin
          valid_240 <= _GEN_4620;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_241 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_241 <= _GEN_2294;
        end else begin
          valid_241 <= _GEN_4621;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_242 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_242 <= _GEN_2295;
        end else begin
          valid_242 <= _GEN_4622;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_243 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_243 <= _GEN_2296;
        end else begin
          valid_243 <= _GEN_4623;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_244 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_244 <= _GEN_2297;
        end else begin
          valid_244 <= _GEN_4624;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_245 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_245 <= _GEN_2298;
        end else begin
          valid_245 <= _GEN_4625;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_246 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_246 <= _GEN_2299;
        end else begin
          valid_246 <= _GEN_4626;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_247 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_247 <= _GEN_2300;
        end else begin
          valid_247 <= _GEN_4627;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_248 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_248 <= _GEN_2301;
        end else begin
          valid_248 <= _GEN_4628;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_249 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_249 <= _GEN_2302;
        end else begin
          valid_249 <= _GEN_4629;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_250 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_250 <= _GEN_2303;
        end else begin
          valid_250 <= _GEN_4630;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_251 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_251 <= _GEN_2304;
        end else begin
          valid_251 <= _GEN_4631;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_252 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_252 <= _GEN_2305;
        end else begin
          valid_252 <= _GEN_4632;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_253 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_253 <= _GEN_2306;
        end else begin
          valid_253 <= _GEN_4633;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_254 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_254 <= _GEN_2307;
        end else begin
          valid_254 <= _GEN_4634;
        end
      end
    end
    if (reset) begin // @[Icache.scala 18:24]
      valid_255 <= 1'h0; // @[Icache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          valid_255 <= _GEN_2308;
        end else begin
          valid_255 <= _GEN_4635;
        end
      end
    end
    if (reset) begin // @[Icache.scala 26:22]
      state <= 3'h0; // @[Icache.scala 26:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_imem_inst_valid) begin // @[Icache.scala 58:28]
        state <= 3'h1; // @[Icache.scala 59:15]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (io_imem_inst_valid) begin // @[Icache.scala 64:28]
        state <= 3'h2; // @[Icache.scala 65:15]
      end else begin
        state <= 3'h0; // @[Icache.scala 68:15]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      state <= _GEN_2052;
    end else begin
      state <= _GEN_4371;
    end
    if (reset) begin // @[Icache.scala 42:28]
      inst_ready <= 1'h0; // @[Icache.scala 42:28]
    end else if (_T) begin // @[Conditional.scala 40:58]
      inst_ready <= 1'h0; // @[Icache.scala 57:18]
    end else if (!(_T_1)) begin // @[Conditional.scala 39:67]
      if (_T_2) begin // @[Conditional.scala 39:67]
        inst_ready <= _GEN_2821;
      end else begin
        inst_ready <= _GEN_4379;
      end
    end
    if (reset) begin // @[Icache.scala 51:28]
      cache_fill <= 1'h0; // @[Icache.scala 51:28]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          cache_fill <= _GEN_4376;
        end
      end
    end
    if (reset) begin // @[Icache.scala 52:28]
      cache_wen <= 1'h0; // @[Icache.scala 52:28]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          cache_wen <= _GEN_4377;
        end
      end
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_wdata <= 128'h0; // @[Icache.scala 53:28]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          cache_wdata <= _GEN_4378;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_0 = _RAND_0[19:0];
  _RAND_1 = {1{`RANDOM}};
  tag_1 = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  tag_2 = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  tag_3 = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  tag_4 = _RAND_4[19:0];
  _RAND_5 = {1{`RANDOM}};
  tag_5 = _RAND_5[19:0];
  _RAND_6 = {1{`RANDOM}};
  tag_6 = _RAND_6[19:0];
  _RAND_7 = {1{`RANDOM}};
  tag_7 = _RAND_7[19:0];
  _RAND_8 = {1{`RANDOM}};
  tag_8 = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  tag_9 = _RAND_9[19:0];
  _RAND_10 = {1{`RANDOM}};
  tag_10 = _RAND_10[19:0];
  _RAND_11 = {1{`RANDOM}};
  tag_11 = _RAND_11[19:0];
  _RAND_12 = {1{`RANDOM}};
  tag_12 = _RAND_12[19:0];
  _RAND_13 = {1{`RANDOM}};
  tag_13 = _RAND_13[19:0];
  _RAND_14 = {1{`RANDOM}};
  tag_14 = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  tag_15 = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  tag_16 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  tag_17 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  tag_18 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  tag_19 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  tag_20 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  tag_21 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  tag_22 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  tag_23 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  tag_24 = _RAND_24[19:0];
  _RAND_25 = {1{`RANDOM}};
  tag_25 = _RAND_25[19:0];
  _RAND_26 = {1{`RANDOM}};
  tag_26 = _RAND_26[19:0];
  _RAND_27 = {1{`RANDOM}};
  tag_27 = _RAND_27[19:0];
  _RAND_28 = {1{`RANDOM}};
  tag_28 = _RAND_28[19:0];
  _RAND_29 = {1{`RANDOM}};
  tag_29 = _RAND_29[19:0];
  _RAND_30 = {1{`RANDOM}};
  tag_30 = _RAND_30[19:0];
  _RAND_31 = {1{`RANDOM}};
  tag_31 = _RAND_31[19:0];
  _RAND_32 = {1{`RANDOM}};
  tag_32 = _RAND_32[19:0];
  _RAND_33 = {1{`RANDOM}};
  tag_33 = _RAND_33[19:0];
  _RAND_34 = {1{`RANDOM}};
  tag_34 = _RAND_34[19:0];
  _RAND_35 = {1{`RANDOM}};
  tag_35 = _RAND_35[19:0];
  _RAND_36 = {1{`RANDOM}};
  tag_36 = _RAND_36[19:0];
  _RAND_37 = {1{`RANDOM}};
  tag_37 = _RAND_37[19:0];
  _RAND_38 = {1{`RANDOM}};
  tag_38 = _RAND_38[19:0];
  _RAND_39 = {1{`RANDOM}};
  tag_39 = _RAND_39[19:0];
  _RAND_40 = {1{`RANDOM}};
  tag_40 = _RAND_40[19:0];
  _RAND_41 = {1{`RANDOM}};
  tag_41 = _RAND_41[19:0];
  _RAND_42 = {1{`RANDOM}};
  tag_42 = _RAND_42[19:0];
  _RAND_43 = {1{`RANDOM}};
  tag_43 = _RAND_43[19:0];
  _RAND_44 = {1{`RANDOM}};
  tag_44 = _RAND_44[19:0];
  _RAND_45 = {1{`RANDOM}};
  tag_45 = _RAND_45[19:0];
  _RAND_46 = {1{`RANDOM}};
  tag_46 = _RAND_46[19:0];
  _RAND_47 = {1{`RANDOM}};
  tag_47 = _RAND_47[19:0];
  _RAND_48 = {1{`RANDOM}};
  tag_48 = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  tag_49 = _RAND_49[19:0];
  _RAND_50 = {1{`RANDOM}};
  tag_50 = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  tag_51 = _RAND_51[19:0];
  _RAND_52 = {1{`RANDOM}};
  tag_52 = _RAND_52[19:0];
  _RAND_53 = {1{`RANDOM}};
  tag_53 = _RAND_53[19:0];
  _RAND_54 = {1{`RANDOM}};
  tag_54 = _RAND_54[19:0];
  _RAND_55 = {1{`RANDOM}};
  tag_55 = _RAND_55[19:0];
  _RAND_56 = {1{`RANDOM}};
  tag_56 = _RAND_56[19:0];
  _RAND_57 = {1{`RANDOM}};
  tag_57 = _RAND_57[19:0];
  _RAND_58 = {1{`RANDOM}};
  tag_58 = _RAND_58[19:0];
  _RAND_59 = {1{`RANDOM}};
  tag_59 = _RAND_59[19:0];
  _RAND_60 = {1{`RANDOM}};
  tag_60 = _RAND_60[19:0];
  _RAND_61 = {1{`RANDOM}};
  tag_61 = _RAND_61[19:0];
  _RAND_62 = {1{`RANDOM}};
  tag_62 = _RAND_62[19:0];
  _RAND_63 = {1{`RANDOM}};
  tag_63 = _RAND_63[19:0];
  _RAND_64 = {1{`RANDOM}};
  tag_64 = _RAND_64[19:0];
  _RAND_65 = {1{`RANDOM}};
  tag_65 = _RAND_65[19:0];
  _RAND_66 = {1{`RANDOM}};
  tag_66 = _RAND_66[19:0];
  _RAND_67 = {1{`RANDOM}};
  tag_67 = _RAND_67[19:0];
  _RAND_68 = {1{`RANDOM}};
  tag_68 = _RAND_68[19:0];
  _RAND_69 = {1{`RANDOM}};
  tag_69 = _RAND_69[19:0];
  _RAND_70 = {1{`RANDOM}};
  tag_70 = _RAND_70[19:0];
  _RAND_71 = {1{`RANDOM}};
  tag_71 = _RAND_71[19:0];
  _RAND_72 = {1{`RANDOM}};
  tag_72 = _RAND_72[19:0];
  _RAND_73 = {1{`RANDOM}};
  tag_73 = _RAND_73[19:0];
  _RAND_74 = {1{`RANDOM}};
  tag_74 = _RAND_74[19:0];
  _RAND_75 = {1{`RANDOM}};
  tag_75 = _RAND_75[19:0];
  _RAND_76 = {1{`RANDOM}};
  tag_76 = _RAND_76[19:0];
  _RAND_77 = {1{`RANDOM}};
  tag_77 = _RAND_77[19:0];
  _RAND_78 = {1{`RANDOM}};
  tag_78 = _RAND_78[19:0];
  _RAND_79 = {1{`RANDOM}};
  tag_79 = _RAND_79[19:0];
  _RAND_80 = {1{`RANDOM}};
  tag_80 = _RAND_80[19:0];
  _RAND_81 = {1{`RANDOM}};
  tag_81 = _RAND_81[19:0];
  _RAND_82 = {1{`RANDOM}};
  tag_82 = _RAND_82[19:0];
  _RAND_83 = {1{`RANDOM}};
  tag_83 = _RAND_83[19:0];
  _RAND_84 = {1{`RANDOM}};
  tag_84 = _RAND_84[19:0];
  _RAND_85 = {1{`RANDOM}};
  tag_85 = _RAND_85[19:0];
  _RAND_86 = {1{`RANDOM}};
  tag_86 = _RAND_86[19:0];
  _RAND_87 = {1{`RANDOM}};
  tag_87 = _RAND_87[19:0];
  _RAND_88 = {1{`RANDOM}};
  tag_88 = _RAND_88[19:0];
  _RAND_89 = {1{`RANDOM}};
  tag_89 = _RAND_89[19:0];
  _RAND_90 = {1{`RANDOM}};
  tag_90 = _RAND_90[19:0];
  _RAND_91 = {1{`RANDOM}};
  tag_91 = _RAND_91[19:0];
  _RAND_92 = {1{`RANDOM}};
  tag_92 = _RAND_92[19:0];
  _RAND_93 = {1{`RANDOM}};
  tag_93 = _RAND_93[19:0];
  _RAND_94 = {1{`RANDOM}};
  tag_94 = _RAND_94[19:0];
  _RAND_95 = {1{`RANDOM}};
  tag_95 = _RAND_95[19:0];
  _RAND_96 = {1{`RANDOM}};
  tag_96 = _RAND_96[19:0];
  _RAND_97 = {1{`RANDOM}};
  tag_97 = _RAND_97[19:0];
  _RAND_98 = {1{`RANDOM}};
  tag_98 = _RAND_98[19:0];
  _RAND_99 = {1{`RANDOM}};
  tag_99 = _RAND_99[19:0];
  _RAND_100 = {1{`RANDOM}};
  tag_100 = _RAND_100[19:0];
  _RAND_101 = {1{`RANDOM}};
  tag_101 = _RAND_101[19:0];
  _RAND_102 = {1{`RANDOM}};
  tag_102 = _RAND_102[19:0];
  _RAND_103 = {1{`RANDOM}};
  tag_103 = _RAND_103[19:0];
  _RAND_104 = {1{`RANDOM}};
  tag_104 = _RAND_104[19:0];
  _RAND_105 = {1{`RANDOM}};
  tag_105 = _RAND_105[19:0];
  _RAND_106 = {1{`RANDOM}};
  tag_106 = _RAND_106[19:0];
  _RAND_107 = {1{`RANDOM}};
  tag_107 = _RAND_107[19:0];
  _RAND_108 = {1{`RANDOM}};
  tag_108 = _RAND_108[19:0];
  _RAND_109 = {1{`RANDOM}};
  tag_109 = _RAND_109[19:0];
  _RAND_110 = {1{`RANDOM}};
  tag_110 = _RAND_110[19:0];
  _RAND_111 = {1{`RANDOM}};
  tag_111 = _RAND_111[19:0];
  _RAND_112 = {1{`RANDOM}};
  tag_112 = _RAND_112[19:0];
  _RAND_113 = {1{`RANDOM}};
  tag_113 = _RAND_113[19:0];
  _RAND_114 = {1{`RANDOM}};
  tag_114 = _RAND_114[19:0];
  _RAND_115 = {1{`RANDOM}};
  tag_115 = _RAND_115[19:0];
  _RAND_116 = {1{`RANDOM}};
  tag_116 = _RAND_116[19:0];
  _RAND_117 = {1{`RANDOM}};
  tag_117 = _RAND_117[19:0];
  _RAND_118 = {1{`RANDOM}};
  tag_118 = _RAND_118[19:0];
  _RAND_119 = {1{`RANDOM}};
  tag_119 = _RAND_119[19:0];
  _RAND_120 = {1{`RANDOM}};
  tag_120 = _RAND_120[19:0];
  _RAND_121 = {1{`RANDOM}};
  tag_121 = _RAND_121[19:0];
  _RAND_122 = {1{`RANDOM}};
  tag_122 = _RAND_122[19:0];
  _RAND_123 = {1{`RANDOM}};
  tag_123 = _RAND_123[19:0];
  _RAND_124 = {1{`RANDOM}};
  tag_124 = _RAND_124[19:0];
  _RAND_125 = {1{`RANDOM}};
  tag_125 = _RAND_125[19:0];
  _RAND_126 = {1{`RANDOM}};
  tag_126 = _RAND_126[19:0];
  _RAND_127 = {1{`RANDOM}};
  tag_127 = _RAND_127[19:0];
  _RAND_128 = {1{`RANDOM}};
  tag_128 = _RAND_128[19:0];
  _RAND_129 = {1{`RANDOM}};
  tag_129 = _RAND_129[19:0];
  _RAND_130 = {1{`RANDOM}};
  tag_130 = _RAND_130[19:0];
  _RAND_131 = {1{`RANDOM}};
  tag_131 = _RAND_131[19:0];
  _RAND_132 = {1{`RANDOM}};
  tag_132 = _RAND_132[19:0];
  _RAND_133 = {1{`RANDOM}};
  tag_133 = _RAND_133[19:0];
  _RAND_134 = {1{`RANDOM}};
  tag_134 = _RAND_134[19:0];
  _RAND_135 = {1{`RANDOM}};
  tag_135 = _RAND_135[19:0];
  _RAND_136 = {1{`RANDOM}};
  tag_136 = _RAND_136[19:0];
  _RAND_137 = {1{`RANDOM}};
  tag_137 = _RAND_137[19:0];
  _RAND_138 = {1{`RANDOM}};
  tag_138 = _RAND_138[19:0];
  _RAND_139 = {1{`RANDOM}};
  tag_139 = _RAND_139[19:0];
  _RAND_140 = {1{`RANDOM}};
  tag_140 = _RAND_140[19:0];
  _RAND_141 = {1{`RANDOM}};
  tag_141 = _RAND_141[19:0];
  _RAND_142 = {1{`RANDOM}};
  tag_142 = _RAND_142[19:0];
  _RAND_143 = {1{`RANDOM}};
  tag_143 = _RAND_143[19:0];
  _RAND_144 = {1{`RANDOM}};
  tag_144 = _RAND_144[19:0];
  _RAND_145 = {1{`RANDOM}};
  tag_145 = _RAND_145[19:0];
  _RAND_146 = {1{`RANDOM}};
  tag_146 = _RAND_146[19:0];
  _RAND_147 = {1{`RANDOM}};
  tag_147 = _RAND_147[19:0];
  _RAND_148 = {1{`RANDOM}};
  tag_148 = _RAND_148[19:0];
  _RAND_149 = {1{`RANDOM}};
  tag_149 = _RAND_149[19:0];
  _RAND_150 = {1{`RANDOM}};
  tag_150 = _RAND_150[19:0];
  _RAND_151 = {1{`RANDOM}};
  tag_151 = _RAND_151[19:0];
  _RAND_152 = {1{`RANDOM}};
  tag_152 = _RAND_152[19:0];
  _RAND_153 = {1{`RANDOM}};
  tag_153 = _RAND_153[19:0];
  _RAND_154 = {1{`RANDOM}};
  tag_154 = _RAND_154[19:0];
  _RAND_155 = {1{`RANDOM}};
  tag_155 = _RAND_155[19:0];
  _RAND_156 = {1{`RANDOM}};
  tag_156 = _RAND_156[19:0];
  _RAND_157 = {1{`RANDOM}};
  tag_157 = _RAND_157[19:0];
  _RAND_158 = {1{`RANDOM}};
  tag_158 = _RAND_158[19:0];
  _RAND_159 = {1{`RANDOM}};
  tag_159 = _RAND_159[19:0];
  _RAND_160 = {1{`RANDOM}};
  tag_160 = _RAND_160[19:0];
  _RAND_161 = {1{`RANDOM}};
  tag_161 = _RAND_161[19:0];
  _RAND_162 = {1{`RANDOM}};
  tag_162 = _RAND_162[19:0];
  _RAND_163 = {1{`RANDOM}};
  tag_163 = _RAND_163[19:0];
  _RAND_164 = {1{`RANDOM}};
  tag_164 = _RAND_164[19:0];
  _RAND_165 = {1{`RANDOM}};
  tag_165 = _RAND_165[19:0];
  _RAND_166 = {1{`RANDOM}};
  tag_166 = _RAND_166[19:0];
  _RAND_167 = {1{`RANDOM}};
  tag_167 = _RAND_167[19:0];
  _RAND_168 = {1{`RANDOM}};
  tag_168 = _RAND_168[19:0];
  _RAND_169 = {1{`RANDOM}};
  tag_169 = _RAND_169[19:0];
  _RAND_170 = {1{`RANDOM}};
  tag_170 = _RAND_170[19:0];
  _RAND_171 = {1{`RANDOM}};
  tag_171 = _RAND_171[19:0];
  _RAND_172 = {1{`RANDOM}};
  tag_172 = _RAND_172[19:0];
  _RAND_173 = {1{`RANDOM}};
  tag_173 = _RAND_173[19:0];
  _RAND_174 = {1{`RANDOM}};
  tag_174 = _RAND_174[19:0];
  _RAND_175 = {1{`RANDOM}};
  tag_175 = _RAND_175[19:0];
  _RAND_176 = {1{`RANDOM}};
  tag_176 = _RAND_176[19:0];
  _RAND_177 = {1{`RANDOM}};
  tag_177 = _RAND_177[19:0];
  _RAND_178 = {1{`RANDOM}};
  tag_178 = _RAND_178[19:0];
  _RAND_179 = {1{`RANDOM}};
  tag_179 = _RAND_179[19:0];
  _RAND_180 = {1{`RANDOM}};
  tag_180 = _RAND_180[19:0];
  _RAND_181 = {1{`RANDOM}};
  tag_181 = _RAND_181[19:0];
  _RAND_182 = {1{`RANDOM}};
  tag_182 = _RAND_182[19:0];
  _RAND_183 = {1{`RANDOM}};
  tag_183 = _RAND_183[19:0];
  _RAND_184 = {1{`RANDOM}};
  tag_184 = _RAND_184[19:0];
  _RAND_185 = {1{`RANDOM}};
  tag_185 = _RAND_185[19:0];
  _RAND_186 = {1{`RANDOM}};
  tag_186 = _RAND_186[19:0];
  _RAND_187 = {1{`RANDOM}};
  tag_187 = _RAND_187[19:0];
  _RAND_188 = {1{`RANDOM}};
  tag_188 = _RAND_188[19:0];
  _RAND_189 = {1{`RANDOM}};
  tag_189 = _RAND_189[19:0];
  _RAND_190 = {1{`RANDOM}};
  tag_190 = _RAND_190[19:0];
  _RAND_191 = {1{`RANDOM}};
  tag_191 = _RAND_191[19:0];
  _RAND_192 = {1{`RANDOM}};
  tag_192 = _RAND_192[19:0];
  _RAND_193 = {1{`RANDOM}};
  tag_193 = _RAND_193[19:0];
  _RAND_194 = {1{`RANDOM}};
  tag_194 = _RAND_194[19:0];
  _RAND_195 = {1{`RANDOM}};
  tag_195 = _RAND_195[19:0];
  _RAND_196 = {1{`RANDOM}};
  tag_196 = _RAND_196[19:0];
  _RAND_197 = {1{`RANDOM}};
  tag_197 = _RAND_197[19:0];
  _RAND_198 = {1{`RANDOM}};
  tag_198 = _RAND_198[19:0];
  _RAND_199 = {1{`RANDOM}};
  tag_199 = _RAND_199[19:0];
  _RAND_200 = {1{`RANDOM}};
  tag_200 = _RAND_200[19:0];
  _RAND_201 = {1{`RANDOM}};
  tag_201 = _RAND_201[19:0];
  _RAND_202 = {1{`RANDOM}};
  tag_202 = _RAND_202[19:0];
  _RAND_203 = {1{`RANDOM}};
  tag_203 = _RAND_203[19:0];
  _RAND_204 = {1{`RANDOM}};
  tag_204 = _RAND_204[19:0];
  _RAND_205 = {1{`RANDOM}};
  tag_205 = _RAND_205[19:0];
  _RAND_206 = {1{`RANDOM}};
  tag_206 = _RAND_206[19:0];
  _RAND_207 = {1{`RANDOM}};
  tag_207 = _RAND_207[19:0];
  _RAND_208 = {1{`RANDOM}};
  tag_208 = _RAND_208[19:0];
  _RAND_209 = {1{`RANDOM}};
  tag_209 = _RAND_209[19:0];
  _RAND_210 = {1{`RANDOM}};
  tag_210 = _RAND_210[19:0];
  _RAND_211 = {1{`RANDOM}};
  tag_211 = _RAND_211[19:0];
  _RAND_212 = {1{`RANDOM}};
  tag_212 = _RAND_212[19:0];
  _RAND_213 = {1{`RANDOM}};
  tag_213 = _RAND_213[19:0];
  _RAND_214 = {1{`RANDOM}};
  tag_214 = _RAND_214[19:0];
  _RAND_215 = {1{`RANDOM}};
  tag_215 = _RAND_215[19:0];
  _RAND_216 = {1{`RANDOM}};
  tag_216 = _RAND_216[19:0];
  _RAND_217 = {1{`RANDOM}};
  tag_217 = _RAND_217[19:0];
  _RAND_218 = {1{`RANDOM}};
  tag_218 = _RAND_218[19:0];
  _RAND_219 = {1{`RANDOM}};
  tag_219 = _RAND_219[19:0];
  _RAND_220 = {1{`RANDOM}};
  tag_220 = _RAND_220[19:0];
  _RAND_221 = {1{`RANDOM}};
  tag_221 = _RAND_221[19:0];
  _RAND_222 = {1{`RANDOM}};
  tag_222 = _RAND_222[19:0];
  _RAND_223 = {1{`RANDOM}};
  tag_223 = _RAND_223[19:0];
  _RAND_224 = {1{`RANDOM}};
  tag_224 = _RAND_224[19:0];
  _RAND_225 = {1{`RANDOM}};
  tag_225 = _RAND_225[19:0];
  _RAND_226 = {1{`RANDOM}};
  tag_226 = _RAND_226[19:0];
  _RAND_227 = {1{`RANDOM}};
  tag_227 = _RAND_227[19:0];
  _RAND_228 = {1{`RANDOM}};
  tag_228 = _RAND_228[19:0];
  _RAND_229 = {1{`RANDOM}};
  tag_229 = _RAND_229[19:0];
  _RAND_230 = {1{`RANDOM}};
  tag_230 = _RAND_230[19:0];
  _RAND_231 = {1{`RANDOM}};
  tag_231 = _RAND_231[19:0];
  _RAND_232 = {1{`RANDOM}};
  tag_232 = _RAND_232[19:0];
  _RAND_233 = {1{`RANDOM}};
  tag_233 = _RAND_233[19:0];
  _RAND_234 = {1{`RANDOM}};
  tag_234 = _RAND_234[19:0];
  _RAND_235 = {1{`RANDOM}};
  tag_235 = _RAND_235[19:0];
  _RAND_236 = {1{`RANDOM}};
  tag_236 = _RAND_236[19:0];
  _RAND_237 = {1{`RANDOM}};
  tag_237 = _RAND_237[19:0];
  _RAND_238 = {1{`RANDOM}};
  tag_238 = _RAND_238[19:0];
  _RAND_239 = {1{`RANDOM}};
  tag_239 = _RAND_239[19:0];
  _RAND_240 = {1{`RANDOM}};
  tag_240 = _RAND_240[19:0];
  _RAND_241 = {1{`RANDOM}};
  tag_241 = _RAND_241[19:0];
  _RAND_242 = {1{`RANDOM}};
  tag_242 = _RAND_242[19:0];
  _RAND_243 = {1{`RANDOM}};
  tag_243 = _RAND_243[19:0];
  _RAND_244 = {1{`RANDOM}};
  tag_244 = _RAND_244[19:0];
  _RAND_245 = {1{`RANDOM}};
  tag_245 = _RAND_245[19:0];
  _RAND_246 = {1{`RANDOM}};
  tag_246 = _RAND_246[19:0];
  _RAND_247 = {1{`RANDOM}};
  tag_247 = _RAND_247[19:0];
  _RAND_248 = {1{`RANDOM}};
  tag_248 = _RAND_248[19:0];
  _RAND_249 = {1{`RANDOM}};
  tag_249 = _RAND_249[19:0];
  _RAND_250 = {1{`RANDOM}};
  tag_250 = _RAND_250[19:0];
  _RAND_251 = {1{`RANDOM}};
  tag_251 = _RAND_251[19:0];
  _RAND_252 = {1{`RANDOM}};
  tag_252 = _RAND_252[19:0];
  _RAND_253 = {1{`RANDOM}};
  tag_253 = _RAND_253[19:0];
  _RAND_254 = {1{`RANDOM}};
  tag_254 = _RAND_254[19:0];
  _RAND_255 = {1{`RANDOM}};
  tag_255 = _RAND_255[19:0];
  _RAND_256 = {1{`RANDOM}};
  valid_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_3 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_4 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_5 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_6 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_7 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_8 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_9 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_10 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_11 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_12 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_13 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_14 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_15 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_16 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_17 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_18 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_19 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_20 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_21 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_22 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_23 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_24 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_25 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_26 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_27 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_28 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_29 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_30 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_31 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_32 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_33 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_34 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_35 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_36 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_37 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_38 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_39 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_40 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_41 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_42 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_43 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_44 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_45 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_46 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_47 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_48 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_49 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_50 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_51 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_52 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_53 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_54 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_55 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_56 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_57 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_58 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_59 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_60 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_61 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_62 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_63 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_64 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_65 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_66 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_67 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid_68 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid_69 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid_70 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid_71 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid_72 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid_73 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid_74 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid_75 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid_76 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid_77 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid_78 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid_79 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid_80 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid_81 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid_82 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid_83 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid_84 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid_85 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid_86 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid_87 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid_88 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid_89 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid_90 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid_91 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid_92 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid_93 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid_94 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid_95 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid_96 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid_97 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid_98 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid_99 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid_100 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid_101 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid_102 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid_103 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid_104 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid_105 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid_106 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid_107 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid_108 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid_109 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid_110 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid_111 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid_112 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid_113 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid_114 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid_115 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid_116 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid_117 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid_118 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid_119 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid_120 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid_121 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid_122 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid_123 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid_124 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid_125 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid_126 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid_127 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  valid_128 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  valid_129 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  valid_130 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  valid_131 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  valid_132 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  valid_133 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  valid_134 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  valid_135 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  valid_136 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  valid_137 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  valid_138 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  valid_139 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  valid_140 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  valid_141 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  valid_142 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  valid_143 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  valid_144 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  valid_145 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  valid_146 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  valid_147 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  valid_148 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  valid_149 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  valid_150 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  valid_151 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  valid_152 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  valid_153 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  valid_154 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  valid_155 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  valid_156 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  valid_157 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  valid_158 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  valid_159 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  valid_160 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  valid_161 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  valid_162 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  valid_163 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  valid_164 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  valid_165 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  valid_166 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  valid_167 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  valid_168 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  valid_169 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  valid_170 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  valid_171 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  valid_172 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  valid_173 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  valid_174 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  valid_175 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  valid_176 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  valid_177 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  valid_178 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  valid_179 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  valid_180 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  valid_181 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  valid_182 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  valid_183 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  valid_184 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  valid_185 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  valid_186 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  valid_187 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  valid_188 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  valid_189 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  valid_190 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  valid_191 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  valid_192 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  valid_193 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  valid_194 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  valid_195 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  valid_196 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  valid_197 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  valid_198 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  valid_199 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  valid_200 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  valid_201 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  valid_202 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  valid_203 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  valid_204 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  valid_205 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  valid_206 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  valid_207 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  valid_208 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  valid_209 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  valid_210 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  valid_211 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  valid_212 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  valid_213 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  valid_214 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  valid_215 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  valid_216 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  valid_217 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  valid_218 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  valid_219 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  valid_220 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  valid_221 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  valid_222 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  valid_223 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  valid_224 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  valid_225 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  valid_226 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  valid_227 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  valid_228 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  valid_229 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  valid_230 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  valid_231 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  valid_232 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  valid_233 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  valid_234 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  valid_235 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  valid_236 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  valid_237 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  valid_238 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  valid_239 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  valid_240 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  valid_241 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  valid_242 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  valid_243 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  valid_244 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  valid_245 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  valid_246 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  valid_247 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  valid_248 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  valid_249 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  valid_250 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  valid_251 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  valid_252 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  valid_253 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  valid_254 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  valid_255 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  state = _RAND_512[2:0];
  _RAND_513 = {1{`RANDOM}};
  inst_ready = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  cache_fill = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  cache_wen = _RAND_515[0:0];
  _RAND_516 = {4{`RANDOM}};
  cache_wdata = _RAND_516[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Dcache(
  input          clock,
  input          reset,
  input          io_dmem_data_valid,
  output         io_dmem_data_ready,
  input          io_dmem_data_req,
  input  [31:0]  io_dmem_data_addr,
  input  [1:0]   io_dmem_data_size,
  input  [7:0]   io_dmem_data_strb,
  output [63:0]  io_dmem_data_read,
  input  [63:0]  io_dmem_data_write,
  output         io_out_data_valid,
  input          io_out_data_ready,
  output         io_out_data_req,
  output [31:0]  io_out_data_addr,
  output [7:0]   io_out_data_strb,
  input  [127:0] io_out_data_read,
  output [127:0] io_out_data_write
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [127:0] _RAND_1028;
  reg [127:0] _RAND_1029;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] req_Q; // @[Dcache.scala 220:19]
  wire  req_CLK; // @[Dcache.scala 220:19]
  wire  req_CEN; // @[Dcache.scala 220:19]
  wire  req_WEN; // @[Dcache.scala 220:19]
  wire [127:0] req_BWEN; // @[Dcache.scala 220:19]
  wire [7:0] req_A; // @[Dcache.scala 220:19]
  wire [127:0] req_D; // @[Dcache.scala 220:19]
  reg [19:0] tag_0; // @[Dcache.scala 16:24]
  reg [19:0] tag_1; // @[Dcache.scala 16:24]
  reg [19:0] tag_2; // @[Dcache.scala 16:24]
  reg [19:0] tag_3; // @[Dcache.scala 16:24]
  reg [19:0] tag_4; // @[Dcache.scala 16:24]
  reg [19:0] tag_5; // @[Dcache.scala 16:24]
  reg [19:0] tag_6; // @[Dcache.scala 16:24]
  reg [19:0] tag_7; // @[Dcache.scala 16:24]
  reg [19:0] tag_8; // @[Dcache.scala 16:24]
  reg [19:0] tag_9; // @[Dcache.scala 16:24]
  reg [19:0] tag_10; // @[Dcache.scala 16:24]
  reg [19:0] tag_11; // @[Dcache.scala 16:24]
  reg [19:0] tag_12; // @[Dcache.scala 16:24]
  reg [19:0] tag_13; // @[Dcache.scala 16:24]
  reg [19:0] tag_14; // @[Dcache.scala 16:24]
  reg [19:0] tag_15; // @[Dcache.scala 16:24]
  reg [19:0] tag_16; // @[Dcache.scala 16:24]
  reg [19:0] tag_17; // @[Dcache.scala 16:24]
  reg [19:0] tag_18; // @[Dcache.scala 16:24]
  reg [19:0] tag_19; // @[Dcache.scala 16:24]
  reg [19:0] tag_20; // @[Dcache.scala 16:24]
  reg [19:0] tag_21; // @[Dcache.scala 16:24]
  reg [19:0] tag_22; // @[Dcache.scala 16:24]
  reg [19:0] tag_23; // @[Dcache.scala 16:24]
  reg [19:0] tag_24; // @[Dcache.scala 16:24]
  reg [19:0] tag_25; // @[Dcache.scala 16:24]
  reg [19:0] tag_26; // @[Dcache.scala 16:24]
  reg [19:0] tag_27; // @[Dcache.scala 16:24]
  reg [19:0] tag_28; // @[Dcache.scala 16:24]
  reg [19:0] tag_29; // @[Dcache.scala 16:24]
  reg [19:0] tag_30; // @[Dcache.scala 16:24]
  reg [19:0] tag_31; // @[Dcache.scala 16:24]
  reg [19:0] tag_32; // @[Dcache.scala 16:24]
  reg [19:0] tag_33; // @[Dcache.scala 16:24]
  reg [19:0] tag_34; // @[Dcache.scala 16:24]
  reg [19:0] tag_35; // @[Dcache.scala 16:24]
  reg [19:0] tag_36; // @[Dcache.scala 16:24]
  reg [19:0] tag_37; // @[Dcache.scala 16:24]
  reg [19:0] tag_38; // @[Dcache.scala 16:24]
  reg [19:0] tag_39; // @[Dcache.scala 16:24]
  reg [19:0] tag_40; // @[Dcache.scala 16:24]
  reg [19:0] tag_41; // @[Dcache.scala 16:24]
  reg [19:0] tag_42; // @[Dcache.scala 16:24]
  reg [19:0] tag_43; // @[Dcache.scala 16:24]
  reg [19:0] tag_44; // @[Dcache.scala 16:24]
  reg [19:0] tag_45; // @[Dcache.scala 16:24]
  reg [19:0] tag_46; // @[Dcache.scala 16:24]
  reg [19:0] tag_47; // @[Dcache.scala 16:24]
  reg [19:0] tag_48; // @[Dcache.scala 16:24]
  reg [19:0] tag_49; // @[Dcache.scala 16:24]
  reg [19:0] tag_50; // @[Dcache.scala 16:24]
  reg [19:0] tag_51; // @[Dcache.scala 16:24]
  reg [19:0] tag_52; // @[Dcache.scala 16:24]
  reg [19:0] tag_53; // @[Dcache.scala 16:24]
  reg [19:0] tag_54; // @[Dcache.scala 16:24]
  reg [19:0] tag_55; // @[Dcache.scala 16:24]
  reg [19:0] tag_56; // @[Dcache.scala 16:24]
  reg [19:0] tag_57; // @[Dcache.scala 16:24]
  reg [19:0] tag_58; // @[Dcache.scala 16:24]
  reg [19:0] tag_59; // @[Dcache.scala 16:24]
  reg [19:0] tag_60; // @[Dcache.scala 16:24]
  reg [19:0] tag_61; // @[Dcache.scala 16:24]
  reg [19:0] tag_62; // @[Dcache.scala 16:24]
  reg [19:0] tag_63; // @[Dcache.scala 16:24]
  reg [19:0] tag_64; // @[Dcache.scala 16:24]
  reg [19:0] tag_65; // @[Dcache.scala 16:24]
  reg [19:0] tag_66; // @[Dcache.scala 16:24]
  reg [19:0] tag_67; // @[Dcache.scala 16:24]
  reg [19:0] tag_68; // @[Dcache.scala 16:24]
  reg [19:0] tag_69; // @[Dcache.scala 16:24]
  reg [19:0] tag_70; // @[Dcache.scala 16:24]
  reg [19:0] tag_71; // @[Dcache.scala 16:24]
  reg [19:0] tag_72; // @[Dcache.scala 16:24]
  reg [19:0] tag_73; // @[Dcache.scala 16:24]
  reg [19:0] tag_74; // @[Dcache.scala 16:24]
  reg [19:0] tag_75; // @[Dcache.scala 16:24]
  reg [19:0] tag_76; // @[Dcache.scala 16:24]
  reg [19:0] tag_77; // @[Dcache.scala 16:24]
  reg [19:0] tag_78; // @[Dcache.scala 16:24]
  reg [19:0] tag_79; // @[Dcache.scala 16:24]
  reg [19:0] tag_80; // @[Dcache.scala 16:24]
  reg [19:0] tag_81; // @[Dcache.scala 16:24]
  reg [19:0] tag_82; // @[Dcache.scala 16:24]
  reg [19:0] tag_83; // @[Dcache.scala 16:24]
  reg [19:0] tag_84; // @[Dcache.scala 16:24]
  reg [19:0] tag_85; // @[Dcache.scala 16:24]
  reg [19:0] tag_86; // @[Dcache.scala 16:24]
  reg [19:0] tag_87; // @[Dcache.scala 16:24]
  reg [19:0] tag_88; // @[Dcache.scala 16:24]
  reg [19:0] tag_89; // @[Dcache.scala 16:24]
  reg [19:0] tag_90; // @[Dcache.scala 16:24]
  reg [19:0] tag_91; // @[Dcache.scala 16:24]
  reg [19:0] tag_92; // @[Dcache.scala 16:24]
  reg [19:0] tag_93; // @[Dcache.scala 16:24]
  reg [19:0] tag_94; // @[Dcache.scala 16:24]
  reg [19:0] tag_95; // @[Dcache.scala 16:24]
  reg [19:0] tag_96; // @[Dcache.scala 16:24]
  reg [19:0] tag_97; // @[Dcache.scala 16:24]
  reg [19:0] tag_98; // @[Dcache.scala 16:24]
  reg [19:0] tag_99; // @[Dcache.scala 16:24]
  reg [19:0] tag_100; // @[Dcache.scala 16:24]
  reg [19:0] tag_101; // @[Dcache.scala 16:24]
  reg [19:0] tag_102; // @[Dcache.scala 16:24]
  reg [19:0] tag_103; // @[Dcache.scala 16:24]
  reg [19:0] tag_104; // @[Dcache.scala 16:24]
  reg [19:0] tag_105; // @[Dcache.scala 16:24]
  reg [19:0] tag_106; // @[Dcache.scala 16:24]
  reg [19:0] tag_107; // @[Dcache.scala 16:24]
  reg [19:0] tag_108; // @[Dcache.scala 16:24]
  reg [19:0] tag_109; // @[Dcache.scala 16:24]
  reg [19:0] tag_110; // @[Dcache.scala 16:24]
  reg [19:0] tag_111; // @[Dcache.scala 16:24]
  reg [19:0] tag_112; // @[Dcache.scala 16:24]
  reg [19:0] tag_113; // @[Dcache.scala 16:24]
  reg [19:0] tag_114; // @[Dcache.scala 16:24]
  reg [19:0] tag_115; // @[Dcache.scala 16:24]
  reg [19:0] tag_116; // @[Dcache.scala 16:24]
  reg [19:0] tag_117; // @[Dcache.scala 16:24]
  reg [19:0] tag_118; // @[Dcache.scala 16:24]
  reg [19:0] tag_119; // @[Dcache.scala 16:24]
  reg [19:0] tag_120; // @[Dcache.scala 16:24]
  reg [19:0] tag_121; // @[Dcache.scala 16:24]
  reg [19:0] tag_122; // @[Dcache.scala 16:24]
  reg [19:0] tag_123; // @[Dcache.scala 16:24]
  reg [19:0] tag_124; // @[Dcache.scala 16:24]
  reg [19:0] tag_125; // @[Dcache.scala 16:24]
  reg [19:0] tag_126; // @[Dcache.scala 16:24]
  reg [19:0] tag_127; // @[Dcache.scala 16:24]
  reg [19:0] tag_128; // @[Dcache.scala 16:24]
  reg [19:0] tag_129; // @[Dcache.scala 16:24]
  reg [19:0] tag_130; // @[Dcache.scala 16:24]
  reg [19:0] tag_131; // @[Dcache.scala 16:24]
  reg [19:0] tag_132; // @[Dcache.scala 16:24]
  reg [19:0] tag_133; // @[Dcache.scala 16:24]
  reg [19:0] tag_134; // @[Dcache.scala 16:24]
  reg [19:0] tag_135; // @[Dcache.scala 16:24]
  reg [19:0] tag_136; // @[Dcache.scala 16:24]
  reg [19:0] tag_137; // @[Dcache.scala 16:24]
  reg [19:0] tag_138; // @[Dcache.scala 16:24]
  reg [19:0] tag_139; // @[Dcache.scala 16:24]
  reg [19:0] tag_140; // @[Dcache.scala 16:24]
  reg [19:0] tag_141; // @[Dcache.scala 16:24]
  reg [19:0] tag_142; // @[Dcache.scala 16:24]
  reg [19:0] tag_143; // @[Dcache.scala 16:24]
  reg [19:0] tag_144; // @[Dcache.scala 16:24]
  reg [19:0] tag_145; // @[Dcache.scala 16:24]
  reg [19:0] tag_146; // @[Dcache.scala 16:24]
  reg [19:0] tag_147; // @[Dcache.scala 16:24]
  reg [19:0] tag_148; // @[Dcache.scala 16:24]
  reg [19:0] tag_149; // @[Dcache.scala 16:24]
  reg [19:0] tag_150; // @[Dcache.scala 16:24]
  reg [19:0] tag_151; // @[Dcache.scala 16:24]
  reg [19:0] tag_152; // @[Dcache.scala 16:24]
  reg [19:0] tag_153; // @[Dcache.scala 16:24]
  reg [19:0] tag_154; // @[Dcache.scala 16:24]
  reg [19:0] tag_155; // @[Dcache.scala 16:24]
  reg [19:0] tag_156; // @[Dcache.scala 16:24]
  reg [19:0] tag_157; // @[Dcache.scala 16:24]
  reg [19:0] tag_158; // @[Dcache.scala 16:24]
  reg [19:0] tag_159; // @[Dcache.scala 16:24]
  reg [19:0] tag_160; // @[Dcache.scala 16:24]
  reg [19:0] tag_161; // @[Dcache.scala 16:24]
  reg [19:0] tag_162; // @[Dcache.scala 16:24]
  reg [19:0] tag_163; // @[Dcache.scala 16:24]
  reg [19:0] tag_164; // @[Dcache.scala 16:24]
  reg [19:0] tag_165; // @[Dcache.scala 16:24]
  reg [19:0] tag_166; // @[Dcache.scala 16:24]
  reg [19:0] tag_167; // @[Dcache.scala 16:24]
  reg [19:0] tag_168; // @[Dcache.scala 16:24]
  reg [19:0] tag_169; // @[Dcache.scala 16:24]
  reg [19:0] tag_170; // @[Dcache.scala 16:24]
  reg [19:0] tag_171; // @[Dcache.scala 16:24]
  reg [19:0] tag_172; // @[Dcache.scala 16:24]
  reg [19:0] tag_173; // @[Dcache.scala 16:24]
  reg [19:0] tag_174; // @[Dcache.scala 16:24]
  reg [19:0] tag_175; // @[Dcache.scala 16:24]
  reg [19:0] tag_176; // @[Dcache.scala 16:24]
  reg [19:0] tag_177; // @[Dcache.scala 16:24]
  reg [19:0] tag_178; // @[Dcache.scala 16:24]
  reg [19:0] tag_179; // @[Dcache.scala 16:24]
  reg [19:0] tag_180; // @[Dcache.scala 16:24]
  reg [19:0] tag_181; // @[Dcache.scala 16:24]
  reg [19:0] tag_182; // @[Dcache.scala 16:24]
  reg [19:0] tag_183; // @[Dcache.scala 16:24]
  reg [19:0] tag_184; // @[Dcache.scala 16:24]
  reg [19:0] tag_185; // @[Dcache.scala 16:24]
  reg [19:0] tag_186; // @[Dcache.scala 16:24]
  reg [19:0] tag_187; // @[Dcache.scala 16:24]
  reg [19:0] tag_188; // @[Dcache.scala 16:24]
  reg [19:0] tag_189; // @[Dcache.scala 16:24]
  reg [19:0] tag_190; // @[Dcache.scala 16:24]
  reg [19:0] tag_191; // @[Dcache.scala 16:24]
  reg [19:0] tag_192; // @[Dcache.scala 16:24]
  reg [19:0] tag_193; // @[Dcache.scala 16:24]
  reg [19:0] tag_194; // @[Dcache.scala 16:24]
  reg [19:0] tag_195; // @[Dcache.scala 16:24]
  reg [19:0] tag_196; // @[Dcache.scala 16:24]
  reg [19:0] tag_197; // @[Dcache.scala 16:24]
  reg [19:0] tag_198; // @[Dcache.scala 16:24]
  reg [19:0] tag_199; // @[Dcache.scala 16:24]
  reg [19:0] tag_200; // @[Dcache.scala 16:24]
  reg [19:0] tag_201; // @[Dcache.scala 16:24]
  reg [19:0] tag_202; // @[Dcache.scala 16:24]
  reg [19:0] tag_203; // @[Dcache.scala 16:24]
  reg [19:0] tag_204; // @[Dcache.scala 16:24]
  reg [19:0] tag_205; // @[Dcache.scala 16:24]
  reg [19:0] tag_206; // @[Dcache.scala 16:24]
  reg [19:0] tag_207; // @[Dcache.scala 16:24]
  reg [19:0] tag_208; // @[Dcache.scala 16:24]
  reg [19:0] tag_209; // @[Dcache.scala 16:24]
  reg [19:0] tag_210; // @[Dcache.scala 16:24]
  reg [19:0] tag_211; // @[Dcache.scala 16:24]
  reg [19:0] tag_212; // @[Dcache.scala 16:24]
  reg [19:0] tag_213; // @[Dcache.scala 16:24]
  reg [19:0] tag_214; // @[Dcache.scala 16:24]
  reg [19:0] tag_215; // @[Dcache.scala 16:24]
  reg [19:0] tag_216; // @[Dcache.scala 16:24]
  reg [19:0] tag_217; // @[Dcache.scala 16:24]
  reg [19:0] tag_218; // @[Dcache.scala 16:24]
  reg [19:0] tag_219; // @[Dcache.scala 16:24]
  reg [19:0] tag_220; // @[Dcache.scala 16:24]
  reg [19:0] tag_221; // @[Dcache.scala 16:24]
  reg [19:0] tag_222; // @[Dcache.scala 16:24]
  reg [19:0] tag_223; // @[Dcache.scala 16:24]
  reg [19:0] tag_224; // @[Dcache.scala 16:24]
  reg [19:0] tag_225; // @[Dcache.scala 16:24]
  reg [19:0] tag_226; // @[Dcache.scala 16:24]
  reg [19:0] tag_227; // @[Dcache.scala 16:24]
  reg [19:0] tag_228; // @[Dcache.scala 16:24]
  reg [19:0] tag_229; // @[Dcache.scala 16:24]
  reg [19:0] tag_230; // @[Dcache.scala 16:24]
  reg [19:0] tag_231; // @[Dcache.scala 16:24]
  reg [19:0] tag_232; // @[Dcache.scala 16:24]
  reg [19:0] tag_233; // @[Dcache.scala 16:24]
  reg [19:0] tag_234; // @[Dcache.scala 16:24]
  reg [19:0] tag_235; // @[Dcache.scala 16:24]
  reg [19:0] tag_236; // @[Dcache.scala 16:24]
  reg [19:0] tag_237; // @[Dcache.scala 16:24]
  reg [19:0] tag_238; // @[Dcache.scala 16:24]
  reg [19:0] tag_239; // @[Dcache.scala 16:24]
  reg [19:0] tag_240; // @[Dcache.scala 16:24]
  reg [19:0] tag_241; // @[Dcache.scala 16:24]
  reg [19:0] tag_242; // @[Dcache.scala 16:24]
  reg [19:0] tag_243; // @[Dcache.scala 16:24]
  reg [19:0] tag_244; // @[Dcache.scala 16:24]
  reg [19:0] tag_245; // @[Dcache.scala 16:24]
  reg [19:0] tag_246; // @[Dcache.scala 16:24]
  reg [19:0] tag_247; // @[Dcache.scala 16:24]
  reg [19:0] tag_248; // @[Dcache.scala 16:24]
  reg [19:0] tag_249; // @[Dcache.scala 16:24]
  reg [19:0] tag_250; // @[Dcache.scala 16:24]
  reg [19:0] tag_251; // @[Dcache.scala 16:24]
  reg [19:0] tag_252; // @[Dcache.scala 16:24]
  reg [19:0] tag_253; // @[Dcache.scala 16:24]
  reg [19:0] tag_254; // @[Dcache.scala 16:24]
  reg [19:0] tag_255; // @[Dcache.scala 16:24]
  reg  valid_0; // @[Dcache.scala 17:24]
  reg  valid_1; // @[Dcache.scala 17:24]
  reg  valid_2; // @[Dcache.scala 17:24]
  reg  valid_3; // @[Dcache.scala 17:24]
  reg  valid_4; // @[Dcache.scala 17:24]
  reg  valid_5; // @[Dcache.scala 17:24]
  reg  valid_6; // @[Dcache.scala 17:24]
  reg  valid_7; // @[Dcache.scala 17:24]
  reg  valid_8; // @[Dcache.scala 17:24]
  reg  valid_9; // @[Dcache.scala 17:24]
  reg  valid_10; // @[Dcache.scala 17:24]
  reg  valid_11; // @[Dcache.scala 17:24]
  reg  valid_12; // @[Dcache.scala 17:24]
  reg  valid_13; // @[Dcache.scala 17:24]
  reg  valid_14; // @[Dcache.scala 17:24]
  reg  valid_15; // @[Dcache.scala 17:24]
  reg  valid_16; // @[Dcache.scala 17:24]
  reg  valid_17; // @[Dcache.scala 17:24]
  reg  valid_18; // @[Dcache.scala 17:24]
  reg  valid_19; // @[Dcache.scala 17:24]
  reg  valid_20; // @[Dcache.scala 17:24]
  reg  valid_21; // @[Dcache.scala 17:24]
  reg  valid_22; // @[Dcache.scala 17:24]
  reg  valid_23; // @[Dcache.scala 17:24]
  reg  valid_24; // @[Dcache.scala 17:24]
  reg  valid_25; // @[Dcache.scala 17:24]
  reg  valid_26; // @[Dcache.scala 17:24]
  reg  valid_27; // @[Dcache.scala 17:24]
  reg  valid_28; // @[Dcache.scala 17:24]
  reg  valid_29; // @[Dcache.scala 17:24]
  reg  valid_30; // @[Dcache.scala 17:24]
  reg  valid_31; // @[Dcache.scala 17:24]
  reg  valid_32; // @[Dcache.scala 17:24]
  reg  valid_33; // @[Dcache.scala 17:24]
  reg  valid_34; // @[Dcache.scala 17:24]
  reg  valid_35; // @[Dcache.scala 17:24]
  reg  valid_36; // @[Dcache.scala 17:24]
  reg  valid_37; // @[Dcache.scala 17:24]
  reg  valid_38; // @[Dcache.scala 17:24]
  reg  valid_39; // @[Dcache.scala 17:24]
  reg  valid_40; // @[Dcache.scala 17:24]
  reg  valid_41; // @[Dcache.scala 17:24]
  reg  valid_42; // @[Dcache.scala 17:24]
  reg  valid_43; // @[Dcache.scala 17:24]
  reg  valid_44; // @[Dcache.scala 17:24]
  reg  valid_45; // @[Dcache.scala 17:24]
  reg  valid_46; // @[Dcache.scala 17:24]
  reg  valid_47; // @[Dcache.scala 17:24]
  reg  valid_48; // @[Dcache.scala 17:24]
  reg  valid_49; // @[Dcache.scala 17:24]
  reg  valid_50; // @[Dcache.scala 17:24]
  reg  valid_51; // @[Dcache.scala 17:24]
  reg  valid_52; // @[Dcache.scala 17:24]
  reg  valid_53; // @[Dcache.scala 17:24]
  reg  valid_54; // @[Dcache.scala 17:24]
  reg  valid_55; // @[Dcache.scala 17:24]
  reg  valid_56; // @[Dcache.scala 17:24]
  reg  valid_57; // @[Dcache.scala 17:24]
  reg  valid_58; // @[Dcache.scala 17:24]
  reg  valid_59; // @[Dcache.scala 17:24]
  reg  valid_60; // @[Dcache.scala 17:24]
  reg  valid_61; // @[Dcache.scala 17:24]
  reg  valid_62; // @[Dcache.scala 17:24]
  reg  valid_63; // @[Dcache.scala 17:24]
  reg  valid_64; // @[Dcache.scala 17:24]
  reg  valid_65; // @[Dcache.scala 17:24]
  reg  valid_66; // @[Dcache.scala 17:24]
  reg  valid_67; // @[Dcache.scala 17:24]
  reg  valid_68; // @[Dcache.scala 17:24]
  reg  valid_69; // @[Dcache.scala 17:24]
  reg  valid_70; // @[Dcache.scala 17:24]
  reg  valid_71; // @[Dcache.scala 17:24]
  reg  valid_72; // @[Dcache.scala 17:24]
  reg  valid_73; // @[Dcache.scala 17:24]
  reg  valid_74; // @[Dcache.scala 17:24]
  reg  valid_75; // @[Dcache.scala 17:24]
  reg  valid_76; // @[Dcache.scala 17:24]
  reg  valid_77; // @[Dcache.scala 17:24]
  reg  valid_78; // @[Dcache.scala 17:24]
  reg  valid_79; // @[Dcache.scala 17:24]
  reg  valid_80; // @[Dcache.scala 17:24]
  reg  valid_81; // @[Dcache.scala 17:24]
  reg  valid_82; // @[Dcache.scala 17:24]
  reg  valid_83; // @[Dcache.scala 17:24]
  reg  valid_84; // @[Dcache.scala 17:24]
  reg  valid_85; // @[Dcache.scala 17:24]
  reg  valid_86; // @[Dcache.scala 17:24]
  reg  valid_87; // @[Dcache.scala 17:24]
  reg  valid_88; // @[Dcache.scala 17:24]
  reg  valid_89; // @[Dcache.scala 17:24]
  reg  valid_90; // @[Dcache.scala 17:24]
  reg  valid_91; // @[Dcache.scala 17:24]
  reg  valid_92; // @[Dcache.scala 17:24]
  reg  valid_93; // @[Dcache.scala 17:24]
  reg  valid_94; // @[Dcache.scala 17:24]
  reg  valid_95; // @[Dcache.scala 17:24]
  reg  valid_96; // @[Dcache.scala 17:24]
  reg  valid_97; // @[Dcache.scala 17:24]
  reg  valid_98; // @[Dcache.scala 17:24]
  reg  valid_99; // @[Dcache.scala 17:24]
  reg  valid_100; // @[Dcache.scala 17:24]
  reg  valid_101; // @[Dcache.scala 17:24]
  reg  valid_102; // @[Dcache.scala 17:24]
  reg  valid_103; // @[Dcache.scala 17:24]
  reg  valid_104; // @[Dcache.scala 17:24]
  reg  valid_105; // @[Dcache.scala 17:24]
  reg  valid_106; // @[Dcache.scala 17:24]
  reg  valid_107; // @[Dcache.scala 17:24]
  reg  valid_108; // @[Dcache.scala 17:24]
  reg  valid_109; // @[Dcache.scala 17:24]
  reg  valid_110; // @[Dcache.scala 17:24]
  reg  valid_111; // @[Dcache.scala 17:24]
  reg  valid_112; // @[Dcache.scala 17:24]
  reg  valid_113; // @[Dcache.scala 17:24]
  reg  valid_114; // @[Dcache.scala 17:24]
  reg  valid_115; // @[Dcache.scala 17:24]
  reg  valid_116; // @[Dcache.scala 17:24]
  reg  valid_117; // @[Dcache.scala 17:24]
  reg  valid_118; // @[Dcache.scala 17:24]
  reg  valid_119; // @[Dcache.scala 17:24]
  reg  valid_120; // @[Dcache.scala 17:24]
  reg  valid_121; // @[Dcache.scala 17:24]
  reg  valid_122; // @[Dcache.scala 17:24]
  reg  valid_123; // @[Dcache.scala 17:24]
  reg  valid_124; // @[Dcache.scala 17:24]
  reg  valid_125; // @[Dcache.scala 17:24]
  reg  valid_126; // @[Dcache.scala 17:24]
  reg  valid_127; // @[Dcache.scala 17:24]
  reg  valid_128; // @[Dcache.scala 17:24]
  reg  valid_129; // @[Dcache.scala 17:24]
  reg  valid_130; // @[Dcache.scala 17:24]
  reg  valid_131; // @[Dcache.scala 17:24]
  reg  valid_132; // @[Dcache.scala 17:24]
  reg  valid_133; // @[Dcache.scala 17:24]
  reg  valid_134; // @[Dcache.scala 17:24]
  reg  valid_135; // @[Dcache.scala 17:24]
  reg  valid_136; // @[Dcache.scala 17:24]
  reg  valid_137; // @[Dcache.scala 17:24]
  reg  valid_138; // @[Dcache.scala 17:24]
  reg  valid_139; // @[Dcache.scala 17:24]
  reg  valid_140; // @[Dcache.scala 17:24]
  reg  valid_141; // @[Dcache.scala 17:24]
  reg  valid_142; // @[Dcache.scala 17:24]
  reg  valid_143; // @[Dcache.scala 17:24]
  reg  valid_144; // @[Dcache.scala 17:24]
  reg  valid_145; // @[Dcache.scala 17:24]
  reg  valid_146; // @[Dcache.scala 17:24]
  reg  valid_147; // @[Dcache.scala 17:24]
  reg  valid_148; // @[Dcache.scala 17:24]
  reg  valid_149; // @[Dcache.scala 17:24]
  reg  valid_150; // @[Dcache.scala 17:24]
  reg  valid_151; // @[Dcache.scala 17:24]
  reg  valid_152; // @[Dcache.scala 17:24]
  reg  valid_153; // @[Dcache.scala 17:24]
  reg  valid_154; // @[Dcache.scala 17:24]
  reg  valid_155; // @[Dcache.scala 17:24]
  reg  valid_156; // @[Dcache.scala 17:24]
  reg  valid_157; // @[Dcache.scala 17:24]
  reg  valid_158; // @[Dcache.scala 17:24]
  reg  valid_159; // @[Dcache.scala 17:24]
  reg  valid_160; // @[Dcache.scala 17:24]
  reg  valid_161; // @[Dcache.scala 17:24]
  reg  valid_162; // @[Dcache.scala 17:24]
  reg  valid_163; // @[Dcache.scala 17:24]
  reg  valid_164; // @[Dcache.scala 17:24]
  reg  valid_165; // @[Dcache.scala 17:24]
  reg  valid_166; // @[Dcache.scala 17:24]
  reg  valid_167; // @[Dcache.scala 17:24]
  reg  valid_168; // @[Dcache.scala 17:24]
  reg  valid_169; // @[Dcache.scala 17:24]
  reg  valid_170; // @[Dcache.scala 17:24]
  reg  valid_171; // @[Dcache.scala 17:24]
  reg  valid_172; // @[Dcache.scala 17:24]
  reg  valid_173; // @[Dcache.scala 17:24]
  reg  valid_174; // @[Dcache.scala 17:24]
  reg  valid_175; // @[Dcache.scala 17:24]
  reg  valid_176; // @[Dcache.scala 17:24]
  reg  valid_177; // @[Dcache.scala 17:24]
  reg  valid_178; // @[Dcache.scala 17:24]
  reg  valid_179; // @[Dcache.scala 17:24]
  reg  valid_180; // @[Dcache.scala 17:24]
  reg  valid_181; // @[Dcache.scala 17:24]
  reg  valid_182; // @[Dcache.scala 17:24]
  reg  valid_183; // @[Dcache.scala 17:24]
  reg  valid_184; // @[Dcache.scala 17:24]
  reg  valid_185; // @[Dcache.scala 17:24]
  reg  valid_186; // @[Dcache.scala 17:24]
  reg  valid_187; // @[Dcache.scala 17:24]
  reg  valid_188; // @[Dcache.scala 17:24]
  reg  valid_189; // @[Dcache.scala 17:24]
  reg  valid_190; // @[Dcache.scala 17:24]
  reg  valid_191; // @[Dcache.scala 17:24]
  reg  valid_192; // @[Dcache.scala 17:24]
  reg  valid_193; // @[Dcache.scala 17:24]
  reg  valid_194; // @[Dcache.scala 17:24]
  reg  valid_195; // @[Dcache.scala 17:24]
  reg  valid_196; // @[Dcache.scala 17:24]
  reg  valid_197; // @[Dcache.scala 17:24]
  reg  valid_198; // @[Dcache.scala 17:24]
  reg  valid_199; // @[Dcache.scala 17:24]
  reg  valid_200; // @[Dcache.scala 17:24]
  reg  valid_201; // @[Dcache.scala 17:24]
  reg  valid_202; // @[Dcache.scala 17:24]
  reg  valid_203; // @[Dcache.scala 17:24]
  reg  valid_204; // @[Dcache.scala 17:24]
  reg  valid_205; // @[Dcache.scala 17:24]
  reg  valid_206; // @[Dcache.scala 17:24]
  reg  valid_207; // @[Dcache.scala 17:24]
  reg  valid_208; // @[Dcache.scala 17:24]
  reg  valid_209; // @[Dcache.scala 17:24]
  reg  valid_210; // @[Dcache.scala 17:24]
  reg  valid_211; // @[Dcache.scala 17:24]
  reg  valid_212; // @[Dcache.scala 17:24]
  reg  valid_213; // @[Dcache.scala 17:24]
  reg  valid_214; // @[Dcache.scala 17:24]
  reg  valid_215; // @[Dcache.scala 17:24]
  reg  valid_216; // @[Dcache.scala 17:24]
  reg  valid_217; // @[Dcache.scala 17:24]
  reg  valid_218; // @[Dcache.scala 17:24]
  reg  valid_219; // @[Dcache.scala 17:24]
  reg  valid_220; // @[Dcache.scala 17:24]
  reg  valid_221; // @[Dcache.scala 17:24]
  reg  valid_222; // @[Dcache.scala 17:24]
  reg  valid_223; // @[Dcache.scala 17:24]
  reg  valid_224; // @[Dcache.scala 17:24]
  reg  valid_225; // @[Dcache.scala 17:24]
  reg  valid_226; // @[Dcache.scala 17:24]
  reg  valid_227; // @[Dcache.scala 17:24]
  reg  valid_228; // @[Dcache.scala 17:24]
  reg  valid_229; // @[Dcache.scala 17:24]
  reg  valid_230; // @[Dcache.scala 17:24]
  reg  valid_231; // @[Dcache.scala 17:24]
  reg  valid_232; // @[Dcache.scala 17:24]
  reg  valid_233; // @[Dcache.scala 17:24]
  reg  valid_234; // @[Dcache.scala 17:24]
  reg  valid_235; // @[Dcache.scala 17:24]
  reg  valid_236; // @[Dcache.scala 17:24]
  reg  valid_237; // @[Dcache.scala 17:24]
  reg  valid_238; // @[Dcache.scala 17:24]
  reg  valid_239; // @[Dcache.scala 17:24]
  reg  valid_240; // @[Dcache.scala 17:24]
  reg  valid_241; // @[Dcache.scala 17:24]
  reg  valid_242; // @[Dcache.scala 17:24]
  reg  valid_243; // @[Dcache.scala 17:24]
  reg  valid_244; // @[Dcache.scala 17:24]
  reg  valid_245; // @[Dcache.scala 17:24]
  reg  valid_246; // @[Dcache.scala 17:24]
  reg  valid_247; // @[Dcache.scala 17:24]
  reg  valid_248; // @[Dcache.scala 17:24]
  reg  valid_249; // @[Dcache.scala 17:24]
  reg  valid_250; // @[Dcache.scala 17:24]
  reg  valid_251; // @[Dcache.scala 17:24]
  reg  valid_252; // @[Dcache.scala 17:24]
  reg  valid_253; // @[Dcache.scala 17:24]
  reg  valid_254; // @[Dcache.scala 17:24]
  reg  valid_255; // @[Dcache.scala 17:24]
  reg  dirty_0; // @[Dcache.scala 18:24]
  reg  dirty_1; // @[Dcache.scala 18:24]
  reg  dirty_2; // @[Dcache.scala 18:24]
  reg  dirty_3; // @[Dcache.scala 18:24]
  reg  dirty_4; // @[Dcache.scala 18:24]
  reg  dirty_5; // @[Dcache.scala 18:24]
  reg  dirty_6; // @[Dcache.scala 18:24]
  reg  dirty_7; // @[Dcache.scala 18:24]
  reg  dirty_8; // @[Dcache.scala 18:24]
  reg  dirty_9; // @[Dcache.scala 18:24]
  reg  dirty_10; // @[Dcache.scala 18:24]
  reg  dirty_11; // @[Dcache.scala 18:24]
  reg  dirty_12; // @[Dcache.scala 18:24]
  reg  dirty_13; // @[Dcache.scala 18:24]
  reg  dirty_14; // @[Dcache.scala 18:24]
  reg  dirty_15; // @[Dcache.scala 18:24]
  reg  dirty_16; // @[Dcache.scala 18:24]
  reg  dirty_17; // @[Dcache.scala 18:24]
  reg  dirty_18; // @[Dcache.scala 18:24]
  reg  dirty_19; // @[Dcache.scala 18:24]
  reg  dirty_20; // @[Dcache.scala 18:24]
  reg  dirty_21; // @[Dcache.scala 18:24]
  reg  dirty_22; // @[Dcache.scala 18:24]
  reg  dirty_23; // @[Dcache.scala 18:24]
  reg  dirty_24; // @[Dcache.scala 18:24]
  reg  dirty_25; // @[Dcache.scala 18:24]
  reg  dirty_26; // @[Dcache.scala 18:24]
  reg  dirty_27; // @[Dcache.scala 18:24]
  reg  dirty_28; // @[Dcache.scala 18:24]
  reg  dirty_29; // @[Dcache.scala 18:24]
  reg  dirty_30; // @[Dcache.scala 18:24]
  reg  dirty_31; // @[Dcache.scala 18:24]
  reg  dirty_32; // @[Dcache.scala 18:24]
  reg  dirty_33; // @[Dcache.scala 18:24]
  reg  dirty_34; // @[Dcache.scala 18:24]
  reg  dirty_35; // @[Dcache.scala 18:24]
  reg  dirty_36; // @[Dcache.scala 18:24]
  reg  dirty_37; // @[Dcache.scala 18:24]
  reg  dirty_38; // @[Dcache.scala 18:24]
  reg  dirty_39; // @[Dcache.scala 18:24]
  reg  dirty_40; // @[Dcache.scala 18:24]
  reg  dirty_41; // @[Dcache.scala 18:24]
  reg  dirty_42; // @[Dcache.scala 18:24]
  reg  dirty_43; // @[Dcache.scala 18:24]
  reg  dirty_44; // @[Dcache.scala 18:24]
  reg  dirty_45; // @[Dcache.scala 18:24]
  reg  dirty_46; // @[Dcache.scala 18:24]
  reg  dirty_47; // @[Dcache.scala 18:24]
  reg  dirty_48; // @[Dcache.scala 18:24]
  reg  dirty_49; // @[Dcache.scala 18:24]
  reg  dirty_50; // @[Dcache.scala 18:24]
  reg  dirty_51; // @[Dcache.scala 18:24]
  reg  dirty_52; // @[Dcache.scala 18:24]
  reg  dirty_53; // @[Dcache.scala 18:24]
  reg  dirty_54; // @[Dcache.scala 18:24]
  reg  dirty_55; // @[Dcache.scala 18:24]
  reg  dirty_56; // @[Dcache.scala 18:24]
  reg  dirty_57; // @[Dcache.scala 18:24]
  reg  dirty_58; // @[Dcache.scala 18:24]
  reg  dirty_59; // @[Dcache.scala 18:24]
  reg  dirty_60; // @[Dcache.scala 18:24]
  reg  dirty_61; // @[Dcache.scala 18:24]
  reg  dirty_62; // @[Dcache.scala 18:24]
  reg  dirty_63; // @[Dcache.scala 18:24]
  reg  dirty_64; // @[Dcache.scala 18:24]
  reg  dirty_65; // @[Dcache.scala 18:24]
  reg  dirty_66; // @[Dcache.scala 18:24]
  reg  dirty_67; // @[Dcache.scala 18:24]
  reg  dirty_68; // @[Dcache.scala 18:24]
  reg  dirty_69; // @[Dcache.scala 18:24]
  reg  dirty_70; // @[Dcache.scala 18:24]
  reg  dirty_71; // @[Dcache.scala 18:24]
  reg  dirty_72; // @[Dcache.scala 18:24]
  reg  dirty_73; // @[Dcache.scala 18:24]
  reg  dirty_74; // @[Dcache.scala 18:24]
  reg  dirty_75; // @[Dcache.scala 18:24]
  reg  dirty_76; // @[Dcache.scala 18:24]
  reg  dirty_77; // @[Dcache.scala 18:24]
  reg  dirty_78; // @[Dcache.scala 18:24]
  reg  dirty_79; // @[Dcache.scala 18:24]
  reg  dirty_80; // @[Dcache.scala 18:24]
  reg  dirty_81; // @[Dcache.scala 18:24]
  reg  dirty_82; // @[Dcache.scala 18:24]
  reg  dirty_83; // @[Dcache.scala 18:24]
  reg  dirty_84; // @[Dcache.scala 18:24]
  reg  dirty_85; // @[Dcache.scala 18:24]
  reg  dirty_86; // @[Dcache.scala 18:24]
  reg  dirty_87; // @[Dcache.scala 18:24]
  reg  dirty_88; // @[Dcache.scala 18:24]
  reg  dirty_89; // @[Dcache.scala 18:24]
  reg  dirty_90; // @[Dcache.scala 18:24]
  reg  dirty_91; // @[Dcache.scala 18:24]
  reg  dirty_92; // @[Dcache.scala 18:24]
  reg  dirty_93; // @[Dcache.scala 18:24]
  reg  dirty_94; // @[Dcache.scala 18:24]
  reg  dirty_95; // @[Dcache.scala 18:24]
  reg  dirty_96; // @[Dcache.scala 18:24]
  reg  dirty_97; // @[Dcache.scala 18:24]
  reg  dirty_98; // @[Dcache.scala 18:24]
  reg  dirty_99; // @[Dcache.scala 18:24]
  reg  dirty_100; // @[Dcache.scala 18:24]
  reg  dirty_101; // @[Dcache.scala 18:24]
  reg  dirty_102; // @[Dcache.scala 18:24]
  reg  dirty_103; // @[Dcache.scala 18:24]
  reg  dirty_104; // @[Dcache.scala 18:24]
  reg  dirty_105; // @[Dcache.scala 18:24]
  reg  dirty_106; // @[Dcache.scala 18:24]
  reg  dirty_107; // @[Dcache.scala 18:24]
  reg  dirty_108; // @[Dcache.scala 18:24]
  reg  dirty_109; // @[Dcache.scala 18:24]
  reg  dirty_110; // @[Dcache.scala 18:24]
  reg  dirty_111; // @[Dcache.scala 18:24]
  reg  dirty_112; // @[Dcache.scala 18:24]
  reg  dirty_113; // @[Dcache.scala 18:24]
  reg  dirty_114; // @[Dcache.scala 18:24]
  reg  dirty_115; // @[Dcache.scala 18:24]
  reg  dirty_116; // @[Dcache.scala 18:24]
  reg  dirty_117; // @[Dcache.scala 18:24]
  reg  dirty_118; // @[Dcache.scala 18:24]
  reg  dirty_119; // @[Dcache.scala 18:24]
  reg  dirty_120; // @[Dcache.scala 18:24]
  reg  dirty_121; // @[Dcache.scala 18:24]
  reg  dirty_122; // @[Dcache.scala 18:24]
  reg  dirty_123; // @[Dcache.scala 18:24]
  reg  dirty_124; // @[Dcache.scala 18:24]
  reg  dirty_125; // @[Dcache.scala 18:24]
  reg  dirty_126; // @[Dcache.scala 18:24]
  reg  dirty_127; // @[Dcache.scala 18:24]
  reg  dirty_128; // @[Dcache.scala 18:24]
  reg  dirty_129; // @[Dcache.scala 18:24]
  reg  dirty_130; // @[Dcache.scala 18:24]
  reg  dirty_131; // @[Dcache.scala 18:24]
  reg  dirty_132; // @[Dcache.scala 18:24]
  reg  dirty_133; // @[Dcache.scala 18:24]
  reg  dirty_134; // @[Dcache.scala 18:24]
  reg  dirty_135; // @[Dcache.scala 18:24]
  reg  dirty_136; // @[Dcache.scala 18:24]
  reg  dirty_137; // @[Dcache.scala 18:24]
  reg  dirty_138; // @[Dcache.scala 18:24]
  reg  dirty_139; // @[Dcache.scala 18:24]
  reg  dirty_140; // @[Dcache.scala 18:24]
  reg  dirty_141; // @[Dcache.scala 18:24]
  reg  dirty_142; // @[Dcache.scala 18:24]
  reg  dirty_143; // @[Dcache.scala 18:24]
  reg  dirty_144; // @[Dcache.scala 18:24]
  reg  dirty_145; // @[Dcache.scala 18:24]
  reg  dirty_146; // @[Dcache.scala 18:24]
  reg  dirty_147; // @[Dcache.scala 18:24]
  reg  dirty_148; // @[Dcache.scala 18:24]
  reg  dirty_149; // @[Dcache.scala 18:24]
  reg  dirty_150; // @[Dcache.scala 18:24]
  reg  dirty_151; // @[Dcache.scala 18:24]
  reg  dirty_152; // @[Dcache.scala 18:24]
  reg  dirty_153; // @[Dcache.scala 18:24]
  reg  dirty_154; // @[Dcache.scala 18:24]
  reg  dirty_155; // @[Dcache.scala 18:24]
  reg  dirty_156; // @[Dcache.scala 18:24]
  reg  dirty_157; // @[Dcache.scala 18:24]
  reg  dirty_158; // @[Dcache.scala 18:24]
  reg  dirty_159; // @[Dcache.scala 18:24]
  reg  dirty_160; // @[Dcache.scala 18:24]
  reg  dirty_161; // @[Dcache.scala 18:24]
  reg  dirty_162; // @[Dcache.scala 18:24]
  reg  dirty_163; // @[Dcache.scala 18:24]
  reg  dirty_164; // @[Dcache.scala 18:24]
  reg  dirty_165; // @[Dcache.scala 18:24]
  reg  dirty_166; // @[Dcache.scala 18:24]
  reg  dirty_167; // @[Dcache.scala 18:24]
  reg  dirty_168; // @[Dcache.scala 18:24]
  reg  dirty_169; // @[Dcache.scala 18:24]
  reg  dirty_170; // @[Dcache.scala 18:24]
  reg  dirty_171; // @[Dcache.scala 18:24]
  reg  dirty_172; // @[Dcache.scala 18:24]
  reg  dirty_173; // @[Dcache.scala 18:24]
  reg  dirty_174; // @[Dcache.scala 18:24]
  reg  dirty_175; // @[Dcache.scala 18:24]
  reg  dirty_176; // @[Dcache.scala 18:24]
  reg  dirty_177; // @[Dcache.scala 18:24]
  reg  dirty_178; // @[Dcache.scala 18:24]
  reg  dirty_179; // @[Dcache.scala 18:24]
  reg  dirty_180; // @[Dcache.scala 18:24]
  reg  dirty_181; // @[Dcache.scala 18:24]
  reg  dirty_182; // @[Dcache.scala 18:24]
  reg  dirty_183; // @[Dcache.scala 18:24]
  reg  dirty_184; // @[Dcache.scala 18:24]
  reg  dirty_185; // @[Dcache.scala 18:24]
  reg  dirty_186; // @[Dcache.scala 18:24]
  reg  dirty_187; // @[Dcache.scala 18:24]
  reg  dirty_188; // @[Dcache.scala 18:24]
  reg  dirty_189; // @[Dcache.scala 18:24]
  reg  dirty_190; // @[Dcache.scala 18:24]
  reg  dirty_191; // @[Dcache.scala 18:24]
  reg  dirty_192; // @[Dcache.scala 18:24]
  reg  dirty_193; // @[Dcache.scala 18:24]
  reg  dirty_194; // @[Dcache.scala 18:24]
  reg  dirty_195; // @[Dcache.scala 18:24]
  reg  dirty_196; // @[Dcache.scala 18:24]
  reg  dirty_197; // @[Dcache.scala 18:24]
  reg  dirty_198; // @[Dcache.scala 18:24]
  reg  dirty_199; // @[Dcache.scala 18:24]
  reg  dirty_200; // @[Dcache.scala 18:24]
  reg  dirty_201; // @[Dcache.scala 18:24]
  reg  dirty_202; // @[Dcache.scala 18:24]
  reg  dirty_203; // @[Dcache.scala 18:24]
  reg  dirty_204; // @[Dcache.scala 18:24]
  reg  dirty_205; // @[Dcache.scala 18:24]
  reg  dirty_206; // @[Dcache.scala 18:24]
  reg  dirty_207; // @[Dcache.scala 18:24]
  reg  dirty_208; // @[Dcache.scala 18:24]
  reg  dirty_209; // @[Dcache.scala 18:24]
  reg  dirty_210; // @[Dcache.scala 18:24]
  reg  dirty_211; // @[Dcache.scala 18:24]
  reg  dirty_212; // @[Dcache.scala 18:24]
  reg  dirty_213; // @[Dcache.scala 18:24]
  reg  dirty_214; // @[Dcache.scala 18:24]
  reg  dirty_215; // @[Dcache.scala 18:24]
  reg  dirty_216; // @[Dcache.scala 18:24]
  reg  dirty_217; // @[Dcache.scala 18:24]
  reg  dirty_218; // @[Dcache.scala 18:24]
  reg  dirty_219; // @[Dcache.scala 18:24]
  reg  dirty_220; // @[Dcache.scala 18:24]
  reg  dirty_221; // @[Dcache.scala 18:24]
  reg  dirty_222; // @[Dcache.scala 18:24]
  reg  dirty_223; // @[Dcache.scala 18:24]
  reg  dirty_224; // @[Dcache.scala 18:24]
  reg  dirty_225; // @[Dcache.scala 18:24]
  reg  dirty_226; // @[Dcache.scala 18:24]
  reg  dirty_227; // @[Dcache.scala 18:24]
  reg  dirty_228; // @[Dcache.scala 18:24]
  reg  dirty_229; // @[Dcache.scala 18:24]
  reg  dirty_230; // @[Dcache.scala 18:24]
  reg  dirty_231; // @[Dcache.scala 18:24]
  reg  dirty_232; // @[Dcache.scala 18:24]
  reg  dirty_233; // @[Dcache.scala 18:24]
  reg  dirty_234; // @[Dcache.scala 18:24]
  reg  dirty_235; // @[Dcache.scala 18:24]
  reg  dirty_236; // @[Dcache.scala 18:24]
  reg  dirty_237; // @[Dcache.scala 18:24]
  reg  dirty_238; // @[Dcache.scala 18:24]
  reg  dirty_239; // @[Dcache.scala 18:24]
  reg  dirty_240; // @[Dcache.scala 18:24]
  reg  dirty_241; // @[Dcache.scala 18:24]
  reg  dirty_242; // @[Dcache.scala 18:24]
  reg  dirty_243; // @[Dcache.scala 18:24]
  reg  dirty_244; // @[Dcache.scala 18:24]
  reg  dirty_245; // @[Dcache.scala 18:24]
  reg  dirty_246; // @[Dcache.scala 18:24]
  reg  dirty_247; // @[Dcache.scala 18:24]
  reg  dirty_248; // @[Dcache.scala 18:24]
  reg  dirty_249; // @[Dcache.scala 18:24]
  reg  dirty_250; // @[Dcache.scala 18:24]
  reg  dirty_251; // @[Dcache.scala 18:24]
  reg  dirty_252; // @[Dcache.scala 18:24]
  reg  dirty_253; // @[Dcache.scala 18:24]
  reg  dirty_254; // @[Dcache.scala 18:24]
  reg  dirty_255; // @[Dcache.scala 18:24]
  reg [3:0] offset_0; // @[Dcache.scala 19:24]
  reg [3:0] offset_1; // @[Dcache.scala 19:24]
  reg [3:0] offset_2; // @[Dcache.scala 19:24]
  reg [3:0] offset_3; // @[Dcache.scala 19:24]
  reg [3:0] offset_4; // @[Dcache.scala 19:24]
  reg [3:0] offset_5; // @[Dcache.scala 19:24]
  reg [3:0] offset_6; // @[Dcache.scala 19:24]
  reg [3:0] offset_7; // @[Dcache.scala 19:24]
  reg [3:0] offset_8; // @[Dcache.scala 19:24]
  reg [3:0] offset_9; // @[Dcache.scala 19:24]
  reg [3:0] offset_10; // @[Dcache.scala 19:24]
  reg [3:0] offset_11; // @[Dcache.scala 19:24]
  reg [3:0] offset_12; // @[Dcache.scala 19:24]
  reg [3:0] offset_13; // @[Dcache.scala 19:24]
  reg [3:0] offset_14; // @[Dcache.scala 19:24]
  reg [3:0] offset_15; // @[Dcache.scala 19:24]
  reg [3:0] offset_16; // @[Dcache.scala 19:24]
  reg [3:0] offset_17; // @[Dcache.scala 19:24]
  reg [3:0] offset_18; // @[Dcache.scala 19:24]
  reg [3:0] offset_19; // @[Dcache.scala 19:24]
  reg [3:0] offset_20; // @[Dcache.scala 19:24]
  reg [3:0] offset_21; // @[Dcache.scala 19:24]
  reg [3:0] offset_22; // @[Dcache.scala 19:24]
  reg [3:0] offset_23; // @[Dcache.scala 19:24]
  reg [3:0] offset_24; // @[Dcache.scala 19:24]
  reg [3:0] offset_25; // @[Dcache.scala 19:24]
  reg [3:0] offset_26; // @[Dcache.scala 19:24]
  reg [3:0] offset_27; // @[Dcache.scala 19:24]
  reg [3:0] offset_28; // @[Dcache.scala 19:24]
  reg [3:0] offset_29; // @[Dcache.scala 19:24]
  reg [3:0] offset_30; // @[Dcache.scala 19:24]
  reg [3:0] offset_31; // @[Dcache.scala 19:24]
  reg [3:0] offset_32; // @[Dcache.scala 19:24]
  reg [3:0] offset_33; // @[Dcache.scala 19:24]
  reg [3:0] offset_34; // @[Dcache.scala 19:24]
  reg [3:0] offset_35; // @[Dcache.scala 19:24]
  reg [3:0] offset_36; // @[Dcache.scala 19:24]
  reg [3:0] offset_37; // @[Dcache.scala 19:24]
  reg [3:0] offset_38; // @[Dcache.scala 19:24]
  reg [3:0] offset_39; // @[Dcache.scala 19:24]
  reg [3:0] offset_40; // @[Dcache.scala 19:24]
  reg [3:0] offset_41; // @[Dcache.scala 19:24]
  reg [3:0] offset_42; // @[Dcache.scala 19:24]
  reg [3:0] offset_43; // @[Dcache.scala 19:24]
  reg [3:0] offset_44; // @[Dcache.scala 19:24]
  reg [3:0] offset_45; // @[Dcache.scala 19:24]
  reg [3:0] offset_46; // @[Dcache.scala 19:24]
  reg [3:0] offset_47; // @[Dcache.scala 19:24]
  reg [3:0] offset_48; // @[Dcache.scala 19:24]
  reg [3:0] offset_49; // @[Dcache.scala 19:24]
  reg [3:0] offset_50; // @[Dcache.scala 19:24]
  reg [3:0] offset_51; // @[Dcache.scala 19:24]
  reg [3:0] offset_52; // @[Dcache.scala 19:24]
  reg [3:0] offset_53; // @[Dcache.scala 19:24]
  reg [3:0] offset_54; // @[Dcache.scala 19:24]
  reg [3:0] offset_55; // @[Dcache.scala 19:24]
  reg [3:0] offset_56; // @[Dcache.scala 19:24]
  reg [3:0] offset_57; // @[Dcache.scala 19:24]
  reg [3:0] offset_58; // @[Dcache.scala 19:24]
  reg [3:0] offset_59; // @[Dcache.scala 19:24]
  reg [3:0] offset_60; // @[Dcache.scala 19:24]
  reg [3:0] offset_61; // @[Dcache.scala 19:24]
  reg [3:0] offset_62; // @[Dcache.scala 19:24]
  reg [3:0] offset_63; // @[Dcache.scala 19:24]
  reg [3:0] offset_64; // @[Dcache.scala 19:24]
  reg [3:0] offset_65; // @[Dcache.scala 19:24]
  reg [3:0] offset_66; // @[Dcache.scala 19:24]
  reg [3:0] offset_67; // @[Dcache.scala 19:24]
  reg [3:0] offset_68; // @[Dcache.scala 19:24]
  reg [3:0] offset_69; // @[Dcache.scala 19:24]
  reg [3:0] offset_70; // @[Dcache.scala 19:24]
  reg [3:0] offset_71; // @[Dcache.scala 19:24]
  reg [3:0] offset_72; // @[Dcache.scala 19:24]
  reg [3:0] offset_73; // @[Dcache.scala 19:24]
  reg [3:0] offset_74; // @[Dcache.scala 19:24]
  reg [3:0] offset_75; // @[Dcache.scala 19:24]
  reg [3:0] offset_76; // @[Dcache.scala 19:24]
  reg [3:0] offset_77; // @[Dcache.scala 19:24]
  reg [3:0] offset_78; // @[Dcache.scala 19:24]
  reg [3:0] offset_79; // @[Dcache.scala 19:24]
  reg [3:0] offset_80; // @[Dcache.scala 19:24]
  reg [3:0] offset_81; // @[Dcache.scala 19:24]
  reg [3:0] offset_82; // @[Dcache.scala 19:24]
  reg [3:0] offset_83; // @[Dcache.scala 19:24]
  reg [3:0] offset_84; // @[Dcache.scala 19:24]
  reg [3:0] offset_85; // @[Dcache.scala 19:24]
  reg [3:0] offset_86; // @[Dcache.scala 19:24]
  reg [3:0] offset_87; // @[Dcache.scala 19:24]
  reg [3:0] offset_88; // @[Dcache.scala 19:24]
  reg [3:0] offset_89; // @[Dcache.scala 19:24]
  reg [3:0] offset_90; // @[Dcache.scala 19:24]
  reg [3:0] offset_91; // @[Dcache.scala 19:24]
  reg [3:0] offset_92; // @[Dcache.scala 19:24]
  reg [3:0] offset_93; // @[Dcache.scala 19:24]
  reg [3:0] offset_94; // @[Dcache.scala 19:24]
  reg [3:0] offset_95; // @[Dcache.scala 19:24]
  reg [3:0] offset_96; // @[Dcache.scala 19:24]
  reg [3:0] offset_97; // @[Dcache.scala 19:24]
  reg [3:0] offset_98; // @[Dcache.scala 19:24]
  reg [3:0] offset_99; // @[Dcache.scala 19:24]
  reg [3:0] offset_100; // @[Dcache.scala 19:24]
  reg [3:0] offset_101; // @[Dcache.scala 19:24]
  reg [3:0] offset_102; // @[Dcache.scala 19:24]
  reg [3:0] offset_103; // @[Dcache.scala 19:24]
  reg [3:0] offset_104; // @[Dcache.scala 19:24]
  reg [3:0] offset_105; // @[Dcache.scala 19:24]
  reg [3:0] offset_106; // @[Dcache.scala 19:24]
  reg [3:0] offset_107; // @[Dcache.scala 19:24]
  reg [3:0] offset_108; // @[Dcache.scala 19:24]
  reg [3:0] offset_109; // @[Dcache.scala 19:24]
  reg [3:0] offset_110; // @[Dcache.scala 19:24]
  reg [3:0] offset_111; // @[Dcache.scala 19:24]
  reg [3:0] offset_112; // @[Dcache.scala 19:24]
  reg [3:0] offset_113; // @[Dcache.scala 19:24]
  reg [3:0] offset_114; // @[Dcache.scala 19:24]
  reg [3:0] offset_115; // @[Dcache.scala 19:24]
  reg [3:0] offset_116; // @[Dcache.scala 19:24]
  reg [3:0] offset_117; // @[Dcache.scala 19:24]
  reg [3:0] offset_118; // @[Dcache.scala 19:24]
  reg [3:0] offset_119; // @[Dcache.scala 19:24]
  reg [3:0] offset_120; // @[Dcache.scala 19:24]
  reg [3:0] offset_121; // @[Dcache.scala 19:24]
  reg [3:0] offset_122; // @[Dcache.scala 19:24]
  reg [3:0] offset_123; // @[Dcache.scala 19:24]
  reg [3:0] offset_124; // @[Dcache.scala 19:24]
  reg [3:0] offset_125; // @[Dcache.scala 19:24]
  reg [3:0] offset_126; // @[Dcache.scala 19:24]
  reg [3:0] offset_127; // @[Dcache.scala 19:24]
  reg [3:0] offset_128; // @[Dcache.scala 19:24]
  reg [3:0] offset_129; // @[Dcache.scala 19:24]
  reg [3:0] offset_130; // @[Dcache.scala 19:24]
  reg [3:0] offset_131; // @[Dcache.scala 19:24]
  reg [3:0] offset_132; // @[Dcache.scala 19:24]
  reg [3:0] offset_133; // @[Dcache.scala 19:24]
  reg [3:0] offset_134; // @[Dcache.scala 19:24]
  reg [3:0] offset_135; // @[Dcache.scala 19:24]
  reg [3:0] offset_136; // @[Dcache.scala 19:24]
  reg [3:0] offset_137; // @[Dcache.scala 19:24]
  reg [3:0] offset_138; // @[Dcache.scala 19:24]
  reg [3:0] offset_139; // @[Dcache.scala 19:24]
  reg [3:0] offset_140; // @[Dcache.scala 19:24]
  reg [3:0] offset_141; // @[Dcache.scala 19:24]
  reg [3:0] offset_142; // @[Dcache.scala 19:24]
  reg [3:0] offset_143; // @[Dcache.scala 19:24]
  reg [3:0] offset_144; // @[Dcache.scala 19:24]
  reg [3:0] offset_145; // @[Dcache.scala 19:24]
  reg [3:0] offset_146; // @[Dcache.scala 19:24]
  reg [3:0] offset_147; // @[Dcache.scala 19:24]
  reg [3:0] offset_148; // @[Dcache.scala 19:24]
  reg [3:0] offset_149; // @[Dcache.scala 19:24]
  reg [3:0] offset_150; // @[Dcache.scala 19:24]
  reg [3:0] offset_151; // @[Dcache.scala 19:24]
  reg [3:0] offset_152; // @[Dcache.scala 19:24]
  reg [3:0] offset_153; // @[Dcache.scala 19:24]
  reg [3:0] offset_154; // @[Dcache.scala 19:24]
  reg [3:0] offset_155; // @[Dcache.scala 19:24]
  reg [3:0] offset_156; // @[Dcache.scala 19:24]
  reg [3:0] offset_157; // @[Dcache.scala 19:24]
  reg [3:0] offset_158; // @[Dcache.scala 19:24]
  reg [3:0] offset_159; // @[Dcache.scala 19:24]
  reg [3:0] offset_160; // @[Dcache.scala 19:24]
  reg [3:0] offset_161; // @[Dcache.scala 19:24]
  reg [3:0] offset_162; // @[Dcache.scala 19:24]
  reg [3:0] offset_163; // @[Dcache.scala 19:24]
  reg [3:0] offset_164; // @[Dcache.scala 19:24]
  reg [3:0] offset_165; // @[Dcache.scala 19:24]
  reg [3:0] offset_166; // @[Dcache.scala 19:24]
  reg [3:0] offset_167; // @[Dcache.scala 19:24]
  reg [3:0] offset_168; // @[Dcache.scala 19:24]
  reg [3:0] offset_169; // @[Dcache.scala 19:24]
  reg [3:0] offset_170; // @[Dcache.scala 19:24]
  reg [3:0] offset_171; // @[Dcache.scala 19:24]
  reg [3:0] offset_172; // @[Dcache.scala 19:24]
  reg [3:0] offset_173; // @[Dcache.scala 19:24]
  reg [3:0] offset_174; // @[Dcache.scala 19:24]
  reg [3:0] offset_175; // @[Dcache.scala 19:24]
  reg [3:0] offset_176; // @[Dcache.scala 19:24]
  reg [3:0] offset_177; // @[Dcache.scala 19:24]
  reg [3:0] offset_178; // @[Dcache.scala 19:24]
  reg [3:0] offset_179; // @[Dcache.scala 19:24]
  reg [3:0] offset_180; // @[Dcache.scala 19:24]
  reg [3:0] offset_181; // @[Dcache.scala 19:24]
  reg [3:0] offset_182; // @[Dcache.scala 19:24]
  reg [3:0] offset_183; // @[Dcache.scala 19:24]
  reg [3:0] offset_184; // @[Dcache.scala 19:24]
  reg [3:0] offset_185; // @[Dcache.scala 19:24]
  reg [3:0] offset_186; // @[Dcache.scala 19:24]
  reg [3:0] offset_187; // @[Dcache.scala 19:24]
  reg [3:0] offset_188; // @[Dcache.scala 19:24]
  reg [3:0] offset_189; // @[Dcache.scala 19:24]
  reg [3:0] offset_190; // @[Dcache.scala 19:24]
  reg [3:0] offset_191; // @[Dcache.scala 19:24]
  reg [3:0] offset_192; // @[Dcache.scala 19:24]
  reg [3:0] offset_193; // @[Dcache.scala 19:24]
  reg [3:0] offset_194; // @[Dcache.scala 19:24]
  reg [3:0] offset_195; // @[Dcache.scala 19:24]
  reg [3:0] offset_196; // @[Dcache.scala 19:24]
  reg [3:0] offset_197; // @[Dcache.scala 19:24]
  reg [3:0] offset_198; // @[Dcache.scala 19:24]
  reg [3:0] offset_199; // @[Dcache.scala 19:24]
  reg [3:0] offset_200; // @[Dcache.scala 19:24]
  reg [3:0] offset_201; // @[Dcache.scala 19:24]
  reg [3:0] offset_202; // @[Dcache.scala 19:24]
  reg [3:0] offset_203; // @[Dcache.scala 19:24]
  reg [3:0] offset_204; // @[Dcache.scala 19:24]
  reg [3:0] offset_205; // @[Dcache.scala 19:24]
  reg [3:0] offset_206; // @[Dcache.scala 19:24]
  reg [3:0] offset_207; // @[Dcache.scala 19:24]
  reg [3:0] offset_208; // @[Dcache.scala 19:24]
  reg [3:0] offset_209; // @[Dcache.scala 19:24]
  reg [3:0] offset_210; // @[Dcache.scala 19:24]
  reg [3:0] offset_211; // @[Dcache.scala 19:24]
  reg [3:0] offset_212; // @[Dcache.scala 19:24]
  reg [3:0] offset_213; // @[Dcache.scala 19:24]
  reg [3:0] offset_214; // @[Dcache.scala 19:24]
  reg [3:0] offset_215; // @[Dcache.scala 19:24]
  reg [3:0] offset_216; // @[Dcache.scala 19:24]
  reg [3:0] offset_217; // @[Dcache.scala 19:24]
  reg [3:0] offset_218; // @[Dcache.scala 19:24]
  reg [3:0] offset_219; // @[Dcache.scala 19:24]
  reg [3:0] offset_220; // @[Dcache.scala 19:24]
  reg [3:0] offset_221; // @[Dcache.scala 19:24]
  reg [3:0] offset_222; // @[Dcache.scala 19:24]
  reg [3:0] offset_223; // @[Dcache.scala 19:24]
  reg [3:0] offset_224; // @[Dcache.scala 19:24]
  reg [3:0] offset_225; // @[Dcache.scala 19:24]
  reg [3:0] offset_226; // @[Dcache.scala 19:24]
  reg [3:0] offset_227; // @[Dcache.scala 19:24]
  reg [3:0] offset_228; // @[Dcache.scala 19:24]
  reg [3:0] offset_229; // @[Dcache.scala 19:24]
  reg [3:0] offset_230; // @[Dcache.scala 19:24]
  reg [3:0] offset_231; // @[Dcache.scala 19:24]
  reg [3:0] offset_232; // @[Dcache.scala 19:24]
  reg [3:0] offset_233; // @[Dcache.scala 19:24]
  reg [3:0] offset_234; // @[Dcache.scala 19:24]
  reg [3:0] offset_235; // @[Dcache.scala 19:24]
  reg [3:0] offset_236; // @[Dcache.scala 19:24]
  reg [3:0] offset_237; // @[Dcache.scala 19:24]
  reg [3:0] offset_238; // @[Dcache.scala 19:24]
  reg [3:0] offset_239; // @[Dcache.scala 19:24]
  reg [3:0] offset_240; // @[Dcache.scala 19:24]
  reg [3:0] offset_241; // @[Dcache.scala 19:24]
  reg [3:0] offset_242; // @[Dcache.scala 19:24]
  reg [3:0] offset_243; // @[Dcache.scala 19:24]
  reg [3:0] offset_244; // @[Dcache.scala 19:24]
  reg [3:0] offset_245; // @[Dcache.scala 19:24]
  reg [3:0] offset_246; // @[Dcache.scala 19:24]
  reg [3:0] offset_247; // @[Dcache.scala 19:24]
  reg [3:0] offset_248; // @[Dcache.scala 19:24]
  reg [3:0] offset_249; // @[Dcache.scala 19:24]
  reg [3:0] offset_250; // @[Dcache.scala 19:24]
  reg [3:0] offset_251; // @[Dcache.scala 19:24]
  reg [3:0] offset_252; // @[Dcache.scala 19:24]
  reg [3:0] offset_253; // @[Dcache.scala 19:24]
  reg [3:0] offset_254; // @[Dcache.scala 19:24]
  reg [3:0] offset_255; // @[Dcache.scala 19:24]
  reg [2:0] state; // @[Dcache.scala 26:22]
  wire [19:0] req_tag = io_dmem_data_addr[31:12]; // @[Dcache.scala 28:30]
  wire [7:0] req_index = io_dmem_data_addr[11:4]; // @[Dcache.scala 29:30]
  wire [3:0] req_offset = io_dmem_data_addr[3:0]; // @[Dcache.scala 30:30]
  wire [19:0] _GEN_1 = 8'h1 == req_index ? tag_1 : tag_0; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_2 = 8'h2 == req_index ? tag_2 : _GEN_1; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_3 = 8'h3 == req_index ? tag_3 : _GEN_2; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_4 = 8'h4 == req_index ? tag_4 : _GEN_3; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_5 = 8'h5 == req_index ? tag_5 : _GEN_4; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_6 = 8'h6 == req_index ? tag_6 : _GEN_5; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_7 = 8'h7 == req_index ? tag_7 : _GEN_6; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_8 = 8'h8 == req_index ? tag_8 : _GEN_7; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_9 = 8'h9 == req_index ? tag_9 : _GEN_8; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_10 = 8'ha == req_index ? tag_10 : _GEN_9; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_11 = 8'hb == req_index ? tag_11 : _GEN_10; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_12 = 8'hc == req_index ? tag_12 : _GEN_11; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_13 = 8'hd == req_index ? tag_13 : _GEN_12; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_14 = 8'he == req_index ? tag_14 : _GEN_13; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_15 = 8'hf == req_index ? tag_15 : _GEN_14; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_16 = 8'h10 == req_index ? tag_16 : _GEN_15; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_17 = 8'h11 == req_index ? tag_17 : _GEN_16; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_18 = 8'h12 == req_index ? tag_18 : _GEN_17; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_19 = 8'h13 == req_index ? tag_19 : _GEN_18; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_20 = 8'h14 == req_index ? tag_20 : _GEN_19; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_21 = 8'h15 == req_index ? tag_21 : _GEN_20; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_22 = 8'h16 == req_index ? tag_22 : _GEN_21; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_23 = 8'h17 == req_index ? tag_23 : _GEN_22; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_24 = 8'h18 == req_index ? tag_24 : _GEN_23; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_25 = 8'h19 == req_index ? tag_25 : _GEN_24; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_26 = 8'h1a == req_index ? tag_26 : _GEN_25; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_27 = 8'h1b == req_index ? tag_27 : _GEN_26; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_28 = 8'h1c == req_index ? tag_28 : _GEN_27; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_29 = 8'h1d == req_index ? tag_29 : _GEN_28; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_30 = 8'h1e == req_index ? tag_30 : _GEN_29; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_31 = 8'h1f == req_index ? tag_31 : _GEN_30; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_32 = 8'h20 == req_index ? tag_32 : _GEN_31; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_33 = 8'h21 == req_index ? tag_33 : _GEN_32; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_34 = 8'h22 == req_index ? tag_34 : _GEN_33; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_35 = 8'h23 == req_index ? tag_35 : _GEN_34; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_36 = 8'h24 == req_index ? tag_36 : _GEN_35; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_37 = 8'h25 == req_index ? tag_37 : _GEN_36; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_38 = 8'h26 == req_index ? tag_38 : _GEN_37; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_39 = 8'h27 == req_index ? tag_39 : _GEN_38; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_40 = 8'h28 == req_index ? tag_40 : _GEN_39; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_41 = 8'h29 == req_index ? tag_41 : _GEN_40; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_42 = 8'h2a == req_index ? tag_42 : _GEN_41; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_43 = 8'h2b == req_index ? tag_43 : _GEN_42; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_44 = 8'h2c == req_index ? tag_44 : _GEN_43; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_45 = 8'h2d == req_index ? tag_45 : _GEN_44; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_46 = 8'h2e == req_index ? tag_46 : _GEN_45; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_47 = 8'h2f == req_index ? tag_47 : _GEN_46; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_48 = 8'h30 == req_index ? tag_48 : _GEN_47; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_49 = 8'h31 == req_index ? tag_49 : _GEN_48; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_50 = 8'h32 == req_index ? tag_50 : _GEN_49; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_51 = 8'h33 == req_index ? tag_51 : _GEN_50; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_52 = 8'h34 == req_index ? tag_52 : _GEN_51; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_53 = 8'h35 == req_index ? tag_53 : _GEN_52; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_54 = 8'h36 == req_index ? tag_54 : _GEN_53; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_55 = 8'h37 == req_index ? tag_55 : _GEN_54; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_56 = 8'h38 == req_index ? tag_56 : _GEN_55; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_57 = 8'h39 == req_index ? tag_57 : _GEN_56; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_58 = 8'h3a == req_index ? tag_58 : _GEN_57; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_59 = 8'h3b == req_index ? tag_59 : _GEN_58; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_60 = 8'h3c == req_index ? tag_60 : _GEN_59; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_61 = 8'h3d == req_index ? tag_61 : _GEN_60; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_62 = 8'h3e == req_index ? tag_62 : _GEN_61; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_63 = 8'h3f == req_index ? tag_63 : _GEN_62; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_64 = 8'h40 == req_index ? tag_64 : _GEN_63; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_65 = 8'h41 == req_index ? tag_65 : _GEN_64; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_66 = 8'h42 == req_index ? tag_66 : _GEN_65; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_67 = 8'h43 == req_index ? tag_67 : _GEN_66; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_68 = 8'h44 == req_index ? tag_68 : _GEN_67; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_69 = 8'h45 == req_index ? tag_69 : _GEN_68; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_70 = 8'h46 == req_index ? tag_70 : _GEN_69; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_71 = 8'h47 == req_index ? tag_71 : _GEN_70; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_72 = 8'h48 == req_index ? tag_72 : _GEN_71; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_73 = 8'h49 == req_index ? tag_73 : _GEN_72; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_74 = 8'h4a == req_index ? tag_74 : _GEN_73; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_75 = 8'h4b == req_index ? tag_75 : _GEN_74; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_76 = 8'h4c == req_index ? tag_76 : _GEN_75; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_77 = 8'h4d == req_index ? tag_77 : _GEN_76; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_78 = 8'h4e == req_index ? tag_78 : _GEN_77; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_79 = 8'h4f == req_index ? tag_79 : _GEN_78; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_80 = 8'h50 == req_index ? tag_80 : _GEN_79; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_81 = 8'h51 == req_index ? tag_81 : _GEN_80; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_82 = 8'h52 == req_index ? tag_82 : _GEN_81; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_83 = 8'h53 == req_index ? tag_83 : _GEN_82; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_84 = 8'h54 == req_index ? tag_84 : _GEN_83; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_85 = 8'h55 == req_index ? tag_85 : _GEN_84; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_86 = 8'h56 == req_index ? tag_86 : _GEN_85; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_87 = 8'h57 == req_index ? tag_87 : _GEN_86; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_88 = 8'h58 == req_index ? tag_88 : _GEN_87; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_89 = 8'h59 == req_index ? tag_89 : _GEN_88; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_90 = 8'h5a == req_index ? tag_90 : _GEN_89; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_91 = 8'h5b == req_index ? tag_91 : _GEN_90; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_92 = 8'h5c == req_index ? tag_92 : _GEN_91; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_93 = 8'h5d == req_index ? tag_93 : _GEN_92; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_94 = 8'h5e == req_index ? tag_94 : _GEN_93; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_95 = 8'h5f == req_index ? tag_95 : _GEN_94; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_96 = 8'h60 == req_index ? tag_96 : _GEN_95; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_97 = 8'h61 == req_index ? tag_97 : _GEN_96; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_98 = 8'h62 == req_index ? tag_98 : _GEN_97; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_99 = 8'h63 == req_index ? tag_99 : _GEN_98; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_100 = 8'h64 == req_index ? tag_100 : _GEN_99; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_101 = 8'h65 == req_index ? tag_101 : _GEN_100; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_102 = 8'h66 == req_index ? tag_102 : _GEN_101; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_103 = 8'h67 == req_index ? tag_103 : _GEN_102; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_104 = 8'h68 == req_index ? tag_104 : _GEN_103; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_105 = 8'h69 == req_index ? tag_105 : _GEN_104; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_106 = 8'h6a == req_index ? tag_106 : _GEN_105; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_107 = 8'h6b == req_index ? tag_107 : _GEN_106; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_108 = 8'h6c == req_index ? tag_108 : _GEN_107; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_109 = 8'h6d == req_index ? tag_109 : _GEN_108; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_110 = 8'h6e == req_index ? tag_110 : _GEN_109; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_111 = 8'h6f == req_index ? tag_111 : _GEN_110; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_112 = 8'h70 == req_index ? tag_112 : _GEN_111; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_113 = 8'h71 == req_index ? tag_113 : _GEN_112; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_114 = 8'h72 == req_index ? tag_114 : _GEN_113; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_115 = 8'h73 == req_index ? tag_115 : _GEN_114; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_116 = 8'h74 == req_index ? tag_116 : _GEN_115; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_117 = 8'h75 == req_index ? tag_117 : _GEN_116; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_118 = 8'h76 == req_index ? tag_118 : _GEN_117; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_119 = 8'h77 == req_index ? tag_119 : _GEN_118; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_120 = 8'h78 == req_index ? tag_120 : _GEN_119; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_121 = 8'h79 == req_index ? tag_121 : _GEN_120; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_122 = 8'h7a == req_index ? tag_122 : _GEN_121; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_123 = 8'h7b == req_index ? tag_123 : _GEN_122; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_124 = 8'h7c == req_index ? tag_124 : _GEN_123; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_125 = 8'h7d == req_index ? tag_125 : _GEN_124; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_126 = 8'h7e == req_index ? tag_126 : _GEN_125; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_127 = 8'h7f == req_index ? tag_127 : _GEN_126; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_128 = 8'h80 == req_index ? tag_128 : _GEN_127; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_129 = 8'h81 == req_index ? tag_129 : _GEN_128; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_130 = 8'h82 == req_index ? tag_130 : _GEN_129; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_131 = 8'h83 == req_index ? tag_131 : _GEN_130; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_132 = 8'h84 == req_index ? tag_132 : _GEN_131; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_133 = 8'h85 == req_index ? tag_133 : _GEN_132; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_134 = 8'h86 == req_index ? tag_134 : _GEN_133; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_135 = 8'h87 == req_index ? tag_135 : _GEN_134; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_136 = 8'h88 == req_index ? tag_136 : _GEN_135; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_137 = 8'h89 == req_index ? tag_137 : _GEN_136; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_138 = 8'h8a == req_index ? tag_138 : _GEN_137; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_139 = 8'h8b == req_index ? tag_139 : _GEN_138; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_140 = 8'h8c == req_index ? tag_140 : _GEN_139; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_141 = 8'h8d == req_index ? tag_141 : _GEN_140; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_142 = 8'h8e == req_index ? tag_142 : _GEN_141; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_143 = 8'h8f == req_index ? tag_143 : _GEN_142; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_144 = 8'h90 == req_index ? tag_144 : _GEN_143; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_145 = 8'h91 == req_index ? tag_145 : _GEN_144; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_146 = 8'h92 == req_index ? tag_146 : _GEN_145; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_147 = 8'h93 == req_index ? tag_147 : _GEN_146; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_148 = 8'h94 == req_index ? tag_148 : _GEN_147; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_149 = 8'h95 == req_index ? tag_149 : _GEN_148; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_150 = 8'h96 == req_index ? tag_150 : _GEN_149; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_151 = 8'h97 == req_index ? tag_151 : _GEN_150; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_152 = 8'h98 == req_index ? tag_152 : _GEN_151; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_153 = 8'h99 == req_index ? tag_153 : _GEN_152; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_154 = 8'h9a == req_index ? tag_154 : _GEN_153; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_155 = 8'h9b == req_index ? tag_155 : _GEN_154; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_156 = 8'h9c == req_index ? tag_156 : _GEN_155; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_157 = 8'h9d == req_index ? tag_157 : _GEN_156; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_158 = 8'h9e == req_index ? tag_158 : _GEN_157; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_159 = 8'h9f == req_index ? tag_159 : _GEN_158; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_160 = 8'ha0 == req_index ? tag_160 : _GEN_159; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_161 = 8'ha1 == req_index ? tag_161 : _GEN_160; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_162 = 8'ha2 == req_index ? tag_162 : _GEN_161; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_163 = 8'ha3 == req_index ? tag_163 : _GEN_162; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_164 = 8'ha4 == req_index ? tag_164 : _GEN_163; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_165 = 8'ha5 == req_index ? tag_165 : _GEN_164; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_166 = 8'ha6 == req_index ? tag_166 : _GEN_165; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_167 = 8'ha7 == req_index ? tag_167 : _GEN_166; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_168 = 8'ha8 == req_index ? tag_168 : _GEN_167; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_169 = 8'ha9 == req_index ? tag_169 : _GEN_168; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_170 = 8'haa == req_index ? tag_170 : _GEN_169; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_171 = 8'hab == req_index ? tag_171 : _GEN_170; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_172 = 8'hac == req_index ? tag_172 : _GEN_171; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_173 = 8'had == req_index ? tag_173 : _GEN_172; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_174 = 8'hae == req_index ? tag_174 : _GEN_173; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_175 = 8'haf == req_index ? tag_175 : _GEN_174; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_176 = 8'hb0 == req_index ? tag_176 : _GEN_175; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_177 = 8'hb1 == req_index ? tag_177 : _GEN_176; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_178 = 8'hb2 == req_index ? tag_178 : _GEN_177; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_179 = 8'hb3 == req_index ? tag_179 : _GEN_178; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_180 = 8'hb4 == req_index ? tag_180 : _GEN_179; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_181 = 8'hb5 == req_index ? tag_181 : _GEN_180; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_182 = 8'hb6 == req_index ? tag_182 : _GEN_181; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_183 = 8'hb7 == req_index ? tag_183 : _GEN_182; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_184 = 8'hb8 == req_index ? tag_184 : _GEN_183; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_185 = 8'hb9 == req_index ? tag_185 : _GEN_184; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_186 = 8'hba == req_index ? tag_186 : _GEN_185; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_187 = 8'hbb == req_index ? tag_187 : _GEN_186; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_188 = 8'hbc == req_index ? tag_188 : _GEN_187; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_189 = 8'hbd == req_index ? tag_189 : _GEN_188; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_190 = 8'hbe == req_index ? tag_190 : _GEN_189; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_191 = 8'hbf == req_index ? tag_191 : _GEN_190; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_192 = 8'hc0 == req_index ? tag_192 : _GEN_191; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_193 = 8'hc1 == req_index ? tag_193 : _GEN_192; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_194 = 8'hc2 == req_index ? tag_194 : _GEN_193; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_195 = 8'hc3 == req_index ? tag_195 : _GEN_194; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_196 = 8'hc4 == req_index ? tag_196 : _GEN_195; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_197 = 8'hc5 == req_index ? tag_197 : _GEN_196; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_198 = 8'hc6 == req_index ? tag_198 : _GEN_197; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_199 = 8'hc7 == req_index ? tag_199 : _GEN_198; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_200 = 8'hc8 == req_index ? tag_200 : _GEN_199; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_201 = 8'hc9 == req_index ? tag_201 : _GEN_200; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_202 = 8'hca == req_index ? tag_202 : _GEN_201; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_203 = 8'hcb == req_index ? tag_203 : _GEN_202; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_204 = 8'hcc == req_index ? tag_204 : _GEN_203; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_205 = 8'hcd == req_index ? tag_205 : _GEN_204; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_206 = 8'hce == req_index ? tag_206 : _GEN_205; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_207 = 8'hcf == req_index ? tag_207 : _GEN_206; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_208 = 8'hd0 == req_index ? tag_208 : _GEN_207; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_209 = 8'hd1 == req_index ? tag_209 : _GEN_208; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_210 = 8'hd2 == req_index ? tag_210 : _GEN_209; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_211 = 8'hd3 == req_index ? tag_211 : _GEN_210; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_212 = 8'hd4 == req_index ? tag_212 : _GEN_211; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_213 = 8'hd5 == req_index ? tag_213 : _GEN_212; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_214 = 8'hd6 == req_index ? tag_214 : _GEN_213; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_215 = 8'hd7 == req_index ? tag_215 : _GEN_214; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_216 = 8'hd8 == req_index ? tag_216 : _GEN_215; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_217 = 8'hd9 == req_index ? tag_217 : _GEN_216; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_218 = 8'hda == req_index ? tag_218 : _GEN_217; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_219 = 8'hdb == req_index ? tag_219 : _GEN_218; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_220 = 8'hdc == req_index ? tag_220 : _GEN_219; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_221 = 8'hdd == req_index ? tag_221 : _GEN_220; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_222 = 8'hde == req_index ? tag_222 : _GEN_221; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_223 = 8'hdf == req_index ? tag_223 : _GEN_222; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_224 = 8'he0 == req_index ? tag_224 : _GEN_223; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_225 = 8'he1 == req_index ? tag_225 : _GEN_224; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_226 = 8'he2 == req_index ? tag_226 : _GEN_225; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_227 = 8'he3 == req_index ? tag_227 : _GEN_226; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_228 = 8'he4 == req_index ? tag_228 : _GEN_227; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_229 = 8'he5 == req_index ? tag_229 : _GEN_228; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_230 = 8'he6 == req_index ? tag_230 : _GEN_229; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_231 = 8'he7 == req_index ? tag_231 : _GEN_230; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_232 = 8'he8 == req_index ? tag_232 : _GEN_231; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_233 = 8'he9 == req_index ? tag_233 : _GEN_232; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_234 = 8'hea == req_index ? tag_234 : _GEN_233; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_235 = 8'heb == req_index ? tag_235 : _GEN_234; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_236 = 8'hec == req_index ? tag_236 : _GEN_235; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_237 = 8'hed == req_index ? tag_237 : _GEN_236; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_238 = 8'hee == req_index ? tag_238 : _GEN_237; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_239 = 8'hef == req_index ? tag_239 : _GEN_238; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_240 = 8'hf0 == req_index ? tag_240 : _GEN_239; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_241 = 8'hf1 == req_index ? tag_241 : _GEN_240; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_242 = 8'hf2 == req_index ? tag_242 : _GEN_241; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_243 = 8'hf3 == req_index ? tag_243 : _GEN_242; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_244 = 8'hf4 == req_index ? tag_244 : _GEN_243; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_245 = 8'hf5 == req_index ? tag_245 : _GEN_244; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_246 = 8'hf6 == req_index ? tag_246 : _GEN_245; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_247 = 8'hf7 == req_index ? tag_247 : _GEN_246; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_248 = 8'hf8 == req_index ? tag_248 : _GEN_247; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_249 = 8'hf9 == req_index ? tag_249 : _GEN_248; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_250 = 8'hfa == req_index ? tag_250 : _GEN_249; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_251 = 8'hfb == req_index ? tag_251 : _GEN_250; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_252 = 8'hfc == req_index ? tag_252 : _GEN_251; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_253 = 8'hfd == req_index ? tag_253 : _GEN_252; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_254 = 8'hfe == req_index ? tag_254 : _GEN_253; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_255 = 8'hff == req_index ? tag_255 : _GEN_254; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire  _GEN_257 = 8'h1 == req_index ? valid_1 : valid_0; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_258 = 8'h2 == req_index ? valid_2 : _GEN_257; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_259 = 8'h3 == req_index ? valid_3 : _GEN_258; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_260 = 8'h4 == req_index ? valid_4 : _GEN_259; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_261 = 8'h5 == req_index ? valid_5 : _GEN_260; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_262 = 8'h6 == req_index ? valid_6 : _GEN_261; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_263 = 8'h7 == req_index ? valid_7 : _GEN_262; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_264 = 8'h8 == req_index ? valid_8 : _GEN_263; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_265 = 8'h9 == req_index ? valid_9 : _GEN_264; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_266 = 8'ha == req_index ? valid_10 : _GEN_265; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_267 = 8'hb == req_index ? valid_11 : _GEN_266; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_268 = 8'hc == req_index ? valid_12 : _GEN_267; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_269 = 8'hd == req_index ? valid_13 : _GEN_268; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_270 = 8'he == req_index ? valid_14 : _GEN_269; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_271 = 8'hf == req_index ? valid_15 : _GEN_270; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_272 = 8'h10 == req_index ? valid_16 : _GEN_271; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_273 = 8'h11 == req_index ? valid_17 : _GEN_272; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_274 = 8'h12 == req_index ? valid_18 : _GEN_273; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_275 = 8'h13 == req_index ? valid_19 : _GEN_274; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_276 = 8'h14 == req_index ? valid_20 : _GEN_275; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_277 = 8'h15 == req_index ? valid_21 : _GEN_276; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_278 = 8'h16 == req_index ? valid_22 : _GEN_277; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_279 = 8'h17 == req_index ? valid_23 : _GEN_278; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_280 = 8'h18 == req_index ? valid_24 : _GEN_279; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_281 = 8'h19 == req_index ? valid_25 : _GEN_280; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_282 = 8'h1a == req_index ? valid_26 : _GEN_281; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_283 = 8'h1b == req_index ? valid_27 : _GEN_282; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_284 = 8'h1c == req_index ? valid_28 : _GEN_283; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_285 = 8'h1d == req_index ? valid_29 : _GEN_284; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_286 = 8'h1e == req_index ? valid_30 : _GEN_285; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_287 = 8'h1f == req_index ? valid_31 : _GEN_286; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_288 = 8'h20 == req_index ? valid_32 : _GEN_287; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_289 = 8'h21 == req_index ? valid_33 : _GEN_288; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_290 = 8'h22 == req_index ? valid_34 : _GEN_289; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_291 = 8'h23 == req_index ? valid_35 : _GEN_290; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_292 = 8'h24 == req_index ? valid_36 : _GEN_291; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_293 = 8'h25 == req_index ? valid_37 : _GEN_292; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_294 = 8'h26 == req_index ? valid_38 : _GEN_293; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_295 = 8'h27 == req_index ? valid_39 : _GEN_294; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_296 = 8'h28 == req_index ? valid_40 : _GEN_295; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_297 = 8'h29 == req_index ? valid_41 : _GEN_296; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_298 = 8'h2a == req_index ? valid_42 : _GEN_297; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_299 = 8'h2b == req_index ? valid_43 : _GEN_298; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_300 = 8'h2c == req_index ? valid_44 : _GEN_299; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_301 = 8'h2d == req_index ? valid_45 : _GEN_300; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_302 = 8'h2e == req_index ? valid_46 : _GEN_301; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_303 = 8'h2f == req_index ? valid_47 : _GEN_302; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_304 = 8'h30 == req_index ? valid_48 : _GEN_303; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_305 = 8'h31 == req_index ? valid_49 : _GEN_304; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_306 = 8'h32 == req_index ? valid_50 : _GEN_305; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_307 = 8'h33 == req_index ? valid_51 : _GEN_306; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_308 = 8'h34 == req_index ? valid_52 : _GEN_307; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_309 = 8'h35 == req_index ? valid_53 : _GEN_308; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_310 = 8'h36 == req_index ? valid_54 : _GEN_309; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_311 = 8'h37 == req_index ? valid_55 : _GEN_310; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_312 = 8'h38 == req_index ? valid_56 : _GEN_311; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_313 = 8'h39 == req_index ? valid_57 : _GEN_312; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_314 = 8'h3a == req_index ? valid_58 : _GEN_313; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_315 = 8'h3b == req_index ? valid_59 : _GEN_314; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_316 = 8'h3c == req_index ? valid_60 : _GEN_315; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_317 = 8'h3d == req_index ? valid_61 : _GEN_316; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_318 = 8'h3e == req_index ? valid_62 : _GEN_317; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_319 = 8'h3f == req_index ? valid_63 : _GEN_318; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_320 = 8'h40 == req_index ? valid_64 : _GEN_319; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_321 = 8'h41 == req_index ? valid_65 : _GEN_320; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_322 = 8'h42 == req_index ? valid_66 : _GEN_321; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_323 = 8'h43 == req_index ? valid_67 : _GEN_322; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_324 = 8'h44 == req_index ? valid_68 : _GEN_323; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_325 = 8'h45 == req_index ? valid_69 : _GEN_324; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_326 = 8'h46 == req_index ? valid_70 : _GEN_325; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_327 = 8'h47 == req_index ? valid_71 : _GEN_326; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_328 = 8'h48 == req_index ? valid_72 : _GEN_327; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_329 = 8'h49 == req_index ? valid_73 : _GEN_328; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_330 = 8'h4a == req_index ? valid_74 : _GEN_329; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_331 = 8'h4b == req_index ? valid_75 : _GEN_330; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_332 = 8'h4c == req_index ? valid_76 : _GEN_331; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_333 = 8'h4d == req_index ? valid_77 : _GEN_332; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_334 = 8'h4e == req_index ? valid_78 : _GEN_333; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_335 = 8'h4f == req_index ? valid_79 : _GEN_334; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_336 = 8'h50 == req_index ? valid_80 : _GEN_335; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_337 = 8'h51 == req_index ? valid_81 : _GEN_336; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_338 = 8'h52 == req_index ? valid_82 : _GEN_337; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_339 = 8'h53 == req_index ? valid_83 : _GEN_338; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_340 = 8'h54 == req_index ? valid_84 : _GEN_339; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_341 = 8'h55 == req_index ? valid_85 : _GEN_340; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_342 = 8'h56 == req_index ? valid_86 : _GEN_341; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_343 = 8'h57 == req_index ? valid_87 : _GEN_342; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_344 = 8'h58 == req_index ? valid_88 : _GEN_343; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_345 = 8'h59 == req_index ? valid_89 : _GEN_344; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_346 = 8'h5a == req_index ? valid_90 : _GEN_345; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_347 = 8'h5b == req_index ? valid_91 : _GEN_346; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_348 = 8'h5c == req_index ? valid_92 : _GEN_347; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_349 = 8'h5d == req_index ? valid_93 : _GEN_348; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_350 = 8'h5e == req_index ? valid_94 : _GEN_349; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_351 = 8'h5f == req_index ? valid_95 : _GEN_350; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_352 = 8'h60 == req_index ? valid_96 : _GEN_351; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_353 = 8'h61 == req_index ? valid_97 : _GEN_352; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_354 = 8'h62 == req_index ? valid_98 : _GEN_353; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_355 = 8'h63 == req_index ? valid_99 : _GEN_354; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_356 = 8'h64 == req_index ? valid_100 : _GEN_355; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_357 = 8'h65 == req_index ? valid_101 : _GEN_356; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_358 = 8'h66 == req_index ? valid_102 : _GEN_357; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_359 = 8'h67 == req_index ? valid_103 : _GEN_358; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_360 = 8'h68 == req_index ? valid_104 : _GEN_359; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_361 = 8'h69 == req_index ? valid_105 : _GEN_360; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_362 = 8'h6a == req_index ? valid_106 : _GEN_361; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_363 = 8'h6b == req_index ? valid_107 : _GEN_362; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_364 = 8'h6c == req_index ? valid_108 : _GEN_363; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_365 = 8'h6d == req_index ? valid_109 : _GEN_364; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_366 = 8'h6e == req_index ? valid_110 : _GEN_365; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_367 = 8'h6f == req_index ? valid_111 : _GEN_366; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_368 = 8'h70 == req_index ? valid_112 : _GEN_367; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_369 = 8'h71 == req_index ? valid_113 : _GEN_368; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_370 = 8'h72 == req_index ? valid_114 : _GEN_369; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_371 = 8'h73 == req_index ? valid_115 : _GEN_370; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_372 = 8'h74 == req_index ? valid_116 : _GEN_371; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_373 = 8'h75 == req_index ? valid_117 : _GEN_372; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_374 = 8'h76 == req_index ? valid_118 : _GEN_373; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_375 = 8'h77 == req_index ? valid_119 : _GEN_374; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_376 = 8'h78 == req_index ? valid_120 : _GEN_375; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_377 = 8'h79 == req_index ? valid_121 : _GEN_376; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_378 = 8'h7a == req_index ? valid_122 : _GEN_377; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_379 = 8'h7b == req_index ? valid_123 : _GEN_378; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_380 = 8'h7c == req_index ? valid_124 : _GEN_379; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_381 = 8'h7d == req_index ? valid_125 : _GEN_380; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_382 = 8'h7e == req_index ? valid_126 : _GEN_381; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_383 = 8'h7f == req_index ? valid_127 : _GEN_382; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_384 = 8'h80 == req_index ? valid_128 : _GEN_383; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_385 = 8'h81 == req_index ? valid_129 : _GEN_384; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_386 = 8'h82 == req_index ? valid_130 : _GEN_385; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_387 = 8'h83 == req_index ? valid_131 : _GEN_386; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_388 = 8'h84 == req_index ? valid_132 : _GEN_387; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_389 = 8'h85 == req_index ? valid_133 : _GEN_388; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_390 = 8'h86 == req_index ? valid_134 : _GEN_389; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_391 = 8'h87 == req_index ? valid_135 : _GEN_390; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_392 = 8'h88 == req_index ? valid_136 : _GEN_391; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_393 = 8'h89 == req_index ? valid_137 : _GEN_392; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_394 = 8'h8a == req_index ? valid_138 : _GEN_393; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_395 = 8'h8b == req_index ? valid_139 : _GEN_394; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_396 = 8'h8c == req_index ? valid_140 : _GEN_395; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_397 = 8'h8d == req_index ? valid_141 : _GEN_396; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_398 = 8'h8e == req_index ? valid_142 : _GEN_397; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_399 = 8'h8f == req_index ? valid_143 : _GEN_398; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_400 = 8'h90 == req_index ? valid_144 : _GEN_399; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_401 = 8'h91 == req_index ? valid_145 : _GEN_400; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_402 = 8'h92 == req_index ? valid_146 : _GEN_401; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_403 = 8'h93 == req_index ? valid_147 : _GEN_402; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_404 = 8'h94 == req_index ? valid_148 : _GEN_403; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_405 = 8'h95 == req_index ? valid_149 : _GEN_404; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_406 = 8'h96 == req_index ? valid_150 : _GEN_405; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_407 = 8'h97 == req_index ? valid_151 : _GEN_406; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_408 = 8'h98 == req_index ? valid_152 : _GEN_407; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_409 = 8'h99 == req_index ? valid_153 : _GEN_408; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_410 = 8'h9a == req_index ? valid_154 : _GEN_409; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_411 = 8'h9b == req_index ? valid_155 : _GEN_410; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_412 = 8'h9c == req_index ? valid_156 : _GEN_411; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_413 = 8'h9d == req_index ? valid_157 : _GEN_412; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_414 = 8'h9e == req_index ? valid_158 : _GEN_413; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_415 = 8'h9f == req_index ? valid_159 : _GEN_414; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_416 = 8'ha0 == req_index ? valid_160 : _GEN_415; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_417 = 8'ha1 == req_index ? valid_161 : _GEN_416; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_418 = 8'ha2 == req_index ? valid_162 : _GEN_417; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_419 = 8'ha3 == req_index ? valid_163 : _GEN_418; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_420 = 8'ha4 == req_index ? valid_164 : _GEN_419; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_421 = 8'ha5 == req_index ? valid_165 : _GEN_420; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_422 = 8'ha6 == req_index ? valid_166 : _GEN_421; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_423 = 8'ha7 == req_index ? valid_167 : _GEN_422; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_424 = 8'ha8 == req_index ? valid_168 : _GEN_423; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_425 = 8'ha9 == req_index ? valid_169 : _GEN_424; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_426 = 8'haa == req_index ? valid_170 : _GEN_425; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_427 = 8'hab == req_index ? valid_171 : _GEN_426; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_428 = 8'hac == req_index ? valid_172 : _GEN_427; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_429 = 8'had == req_index ? valid_173 : _GEN_428; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_430 = 8'hae == req_index ? valid_174 : _GEN_429; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_431 = 8'haf == req_index ? valid_175 : _GEN_430; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_432 = 8'hb0 == req_index ? valid_176 : _GEN_431; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_433 = 8'hb1 == req_index ? valid_177 : _GEN_432; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_434 = 8'hb2 == req_index ? valid_178 : _GEN_433; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_435 = 8'hb3 == req_index ? valid_179 : _GEN_434; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_436 = 8'hb4 == req_index ? valid_180 : _GEN_435; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_437 = 8'hb5 == req_index ? valid_181 : _GEN_436; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_438 = 8'hb6 == req_index ? valid_182 : _GEN_437; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_439 = 8'hb7 == req_index ? valid_183 : _GEN_438; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_440 = 8'hb8 == req_index ? valid_184 : _GEN_439; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_441 = 8'hb9 == req_index ? valid_185 : _GEN_440; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_442 = 8'hba == req_index ? valid_186 : _GEN_441; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_443 = 8'hbb == req_index ? valid_187 : _GEN_442; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_444 = 8'hbc == req_index ? valid_188 : _GEN_443; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_445 = 8'hbd == req_index ? valid_189 : _GEN_444; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_446 = 8'hbe == req_index ? valid_190 : _GEN_445; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_447 = 8'hbf == req_index ? valid_191 : _GEN_446; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_448 = 8'hc0 == req_index ? valid_192 : _GEN_447; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_449 = 8'hc1 == req_index ? valid_193 : _GEN_448; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_450 = 8'hc2 == req_index ? valid_194 : _GEN_449; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_451 = 8'hc3 == req_index ? valid_195 : _GEN_450; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_452 = 8'hc4 == req_index ? valid_196 : _GEN_451; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_453 = 8'hc5 == req_index ? valid_197 : _GEN_452; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_454 = 8'hc6 == req_index ? valid_198 : _GEN_453; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_455 = 8'hc7 == req_index ? valid_199 : _GEN_454; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_456 = 8'hc8 == req_index ? valid_200 : _GEN_455; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_457 = 8'hc9 == req_index ? valid_201 : _GEN_456; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_458 = 8'hca == req_index ? valid_202 : _GEN_457; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_459 = 8'hcb == req_index ? valid_203 : _GEN_458; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_460 = 8'hcc == req_index ? valid_204 : _GEN_459; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_461 = 8'hcd == req_index ? valid_205 : _GEN_460; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_462 = 8'hce == req_index ? valid_206 : _GEN_461; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_463 = 8'hcf == req_index ? valid_207 : _GEN_462; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_464 = 8'hd0 == req_index ? valid_208 : _GEN_463; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_465 = 8'hd1 == req_index ? valid_209 : _GEN_464; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_466 = 8'hd2 == req_index ? valid_210 : _GEN_465; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_467 = 8'hd3 == req_index ? valid_211 : _GEN_466; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_468 = 8'hd4 == req_index ? valid_212 : _GEN_467; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_469 = 8'hd5 == req_index ? valid_213 : _GEN_468; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_470 = 8'hd6 == req_index ? valid_214 : _GEN_469; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_471 = 8'hd7 == req_index ? valid_215 : _GEN_470; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_472 = 8'hd8 == req_index ? valid_216 : _GEN_471; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_473 = 8'hd9 == req_index ? valid_217 : _GEN_472; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_474 = 8'hda == req_index ? valid_218 : _GEN_473; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_475 = 8'hdb == req_index ? valid_219 : _GEN_474; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_476 = 8'hdc == req_index ? valid_220 : _GEN_475; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_477 = 8'hdd == req_index ? valid_221 : _GEN_476; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_478 = 8'hde == req_index ? valid_222 : _GEN_477; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_479 = 8'hdf == req_index ? valid_223 : _GEN_478; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_480 = 8'he0 == req_index ? valid_224 : _GEN_479; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_481 = 8'he1 == req_index ? valid_225 : _GEN_480; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_482 = 8'he2 == req_index ? valid_226 : _GEN_481; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_483 = 8'he3 == req_index ? valid_227 : _GEN_482; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_484 = 8'he4 == req_index ? valid_228 : _GEN_483; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_485 = 8'he5 == req_index ? valid_229 : _GEN_484; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_486 = 8'he6 == req_index ? valid_230 : _GEN_485; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_487 = 8'he7 == req_index ? valid_231 : _GEN_486; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_488 = 8'he8 == req_index ? valid_232 : _GEN_487; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_489 = 8'he9 == req_index ? valid_233 : _GEN_488; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_490 = 8'hea == req_index ? valid_234 : _GEN_489; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_491 = 8'heb == req_index ? valid_235 : _GEN_490; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_492 = 8'hec == req_index ? valid_236 : _GEN_491; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_493 = 8'hed == req_index ? valid_237 : _GEN_492; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_494 = 8'hee == req_index ? valid_238 : _GEN_493; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_495 = 8'hef == req_index ? valid_239 : _GEN_494; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_496 = 8'hf0 == req_index ? valid_240 : _GEN_495; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_497 = 8'hf1 == req_index ? valid_241 : _GEN_496; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_498 = 8'hf2 == req_index ? valid_242 : _GEN_497; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_499 = 8'hf3 == req_index ? valid_243 : _GEN_498; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_500 = 8'hf4 == req_index ? valid_244 : _GEN_499; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_501 = 8'hf5 == req_index ? valid_245 : _GEN_500; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_502 = 8'hf6 == req_index ? valid_246 : _GEN_501; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_503 = 8'hf7 == req_index ? valid_247 : _GEN_502; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_504 = 8'hf8 == req_index ? valid_248 : _GEN_503; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_505 = 8'hf9 == req_index ? valid_249 : _GEN_504; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_506 = 8'hfa == req_index ? valid_250 : _GEN_505; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_507 = 8'hfb == req_index ? valid_251 : _GEN_506; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_508 = 8'hfc == req_index ? valid_252 : _GEN_507; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_509 = 8'hfd == req_index ? valid_253 : _GEN_508; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_510 = 8'hfe == req_index ? valid_254 : _GEN_509; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_511 = 8'hff == req_index ? valid_255 : _GEN_510; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _cache_hit_T_2 = state == 3'h1; // @[Dcache.scala 34:78]
  wire  cache_hit = _GEN_255 == req_tag & _GEN_511 & state == 3'h1; // @[Dcache.scala 34:69]
  wire  _GEN_513 = 8'h1 == req_index ? dirty_1 : dirty_0; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_514 = 8'h2 == req_index ? dirty_2 : _GEN_513; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_515 = 8'h3 == req_index ? dirty_3 : _GEN_514; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_516 = 8'h4 == req_index ? dirty_4 : _GEN_515; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_517 = 8'h5 == req_index ? dirty_5 : _GEN_516; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_518 = 8'h6 == req_index ? dirty_6 : _GEN_517; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_519 = 8'h7 == req_index ? dirty_7 : _GEN_518; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_520 = 8'h8 == req_index ? dirty_8 : _GEN_519; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_521 = 8'h9 == req_index ? dirty_9 : _GEN_520; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_522 = 8'ha == req_index ? dirty_10 : _GEN_521; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_523 = 8'hb == req_index ? dirty_11 : _GEN_522; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_524 = 8'hc == req_index ? dirty_12 : _GEN_523; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_525 = 8'hd == req_index ? dirty_13 : _GEN_524; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_526 = 8'he == req_index ? dirty_14 : _GEN_525; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_527 = 8'hf == req_index ? dirty_15 : _GEN_526; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_528 = 8'h10 == req_index ? dirty_16 : _GEN_527; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_529 = 8'h11 == req_index ? dirty_17 : _GEN_528; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_530 = 8'h12 == req_index ? dirty_18 : _GEN_529; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_531 = 8'h13 == req_index ? dirty_19 : _GEN_530; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_532 = 8'h14 == req_index ? dirty_20 : _GEN_531; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_533 = 8'h15 == req_index ? dirty_21 : _GEN_532; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_534 = 8'h16 == req_index ? dirty_22 : _GEN_533; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_535 = 8'h17 == req_index ? dirty_23 : _GEN_534; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_536 = 8'h18 == req_index ? dirty_24 : _GEN_535; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_537 = 8'h19 == req_index ? dirty_25 : _GEN_536; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_538 = 8'h1a == req_index ? dirty_26 : _GEN_537; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_539 = 8'h1b == req_index ? dirty_27 : _GEN_538; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_540 = 8'h1c == req_index ? dirty_28 : _GEN_539; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_541 = 8'h1d == req_index ? dirty_29 : _GEN_540; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_542 = 8'h1e == req_index ? dirty_30 : _GEN_541; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_543 = 8'h1f == req_index ? dirty_31 : _GEN_542; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_544 = 8'h20 == req_index ? dirty_32 : _GEN_543; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_545 = 8'h21 == req_index ? dirty_33 : _GEN_544; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_546 = 8'h22 == req_index ? dirty_34 : _GEN_545; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_547 = 8'h23 == req_index ? dirty_35 : _GEN_546; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_548 = 8'h24 == req_index ? dirty_36 : _GEN_547; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_549 = 8'h25 == req_index ? dirty_37 : _GEN_548; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_550 = 8'h26 == req_index ? dirty_38 : _GEN_549; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_551 = 8'h27 == req_index ? dirty_39 : _GEN_550; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_552 = 8'h28 == req_index ? dirty_40 : _GEN_551; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_553 = 8'h29 == req_index ? dirty_41 : _GEN_552; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_554 = 8'h2a == req_index ? dirty_42 : _GEN_553; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_555 = 8'h2b == req_index ? dirty_43 : _GEN_554; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_556 = 8'h2c == req_index ? dirty_44 : _GEN_555; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_557 = 8'h2d == req_index ? dirty_45 : _GEN_556; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_558 = 8'h2e == req_index ? dirty_46 : _GEN_557; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_559 = 8'h2f == req_index ? dirty_47 : _GEN_558; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_560 = 8'h30 == req_index ? dirty_48 : _GEN_559; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_561 = 8'h31 == req_index ? dirty_49 : _GEN_560; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_562 = 8'h32 == req_index ? dirty_50 : _GEN_561; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_563 = 8'h33 == req_index ? dirty_51 : _GEN_562; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_564 = 8'h34 == req_index ? dirty_52 : _GEN_563; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_565 = 8'h35 == req_index ? dirty_53 : _GEN_564; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_566 = 8'h36 == req_index ? dirty_54 : _GEN_565; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_567 = 8'h37 == req_index ? dirty_55 : _GEN_566; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_568 = 8'h38 == req_index ? dirty_56 : _GEN_567; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_569 = 8'h39 == req_index ? dirty_57 : _GEN_568; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_570 = 8'h3a == req_index ? dirty_58 : _GEN_569; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_571 = 8'h3b == req_index ? dirty_59 : _GEN_570; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_572 = 8'h3c == req_index ? dirty_60 : _GEN_571; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_573 = 8'h3d == req_index ? dirty_61 : _GEN_572; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_574 = 8'h3e == req_index ? dirty_62 : _GEN_573; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_575 = 8'h3f == req_index ? dirty_63 : _GEN_574; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_576 = 8'h40 == req_index ? dirty_64 : _GEN_575; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_577 = 8'h41 == req_index ? dirty_65 : _GEN_576; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_578 = 8'h42 == req_index ? dirty_66 : _GEN_577; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_579 = 8'h43 == req_index ? dirty_67 : _GEN_578; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_580 = 8'h44 == req_index ? dirty_68 : _GEN_579; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_581 = 8'h45 == req_index ? dirty_69 : _GEN_580; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_582 = 8'h46 == req_index ? dirty_70 : _GEN_581; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_583 = 8'h47 == req_index ? dirty_71 : _GEN_582; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_584 = 8'h48 == req_index ? dirty_72 : _GEN_583; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_585 = 8'h49 == req_index ? dirty_73 : _GEN_584; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_586 = 8'h4a == req_index ? dirty_74 : _GEN_585; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_587 = 8'h4b == req_index ? dirty_75 : _GEN_586; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_588 = 8'h4c == req_index ? dirty_76 : _GEN_587; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_589 = 8'h4d == req_index ? dirty_77 : _GEN_588; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_590 = 8'h4e == req_index ? dirty_78 : _GEN_589; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_591 = 8'h4f == req_index ? dirty_79 : _GEN_590; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_592 = 8'h50 == req_index ? dirty_80 : _GEN_591; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_593 = 8'h51 == req_index ? dirty_81 : _GEN_592; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_594 = 8'h52 == req_index ? dirty_82 : _GEN_593; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_595 = 8'h53 == req_index ? dirty_83 : _GEN_594; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_596 = 8'h54 == req_index ? dirty_84 : _GEN_595; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_597 = 8'h55 == req_index ? dirty_85 : _GEN_596; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_598 = 8'h56 == req_index ? dirty_86 : _GEN_597; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_599 = 8'h57 == req_index ? dirty_87 : _GEN_598; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_600 = 8'h58 == req_index ? dirty_88 : _GEN_599; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_601 = 8'h59 == req_index ? dirty_89 : _GEN_600; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_602 = 8'h5a == req_index ? dirty_90 : _GEN_601; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_603 = 8'h5b == req_index ? dirty_91 : _GEN_602; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_604 = 8'h5c == req_index ? dirty_92 : _GEN_603; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_605 = 8'h5d == req_index ? dirty_93 : _GEN_604; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_606 = 8'h5e == req_index ? dirty_94 : _GEN_605; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_607 = 8'h5f == req_index ? dirty_95 : _GEN_606; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_608 = 8'h60 == req_index ? dirty_96 : _GEN_607; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_609 = 8'h61 == req_index ? dirty_97 : _GEN_608; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_610 = 8'h62 == req_index ? dirty_98 : _GEN_609; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_611 = 8'h63 == req_index ? dirty_99 : _GEN_610; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_612 = 8'h64 == req_index ? dirty_100 : _GEN_611; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_613 = 8'h65 == req_index ? dirty_101 : _GEN_612; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_614 = 8'h66 == req_index ? dirty_102 : _GEN_613; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_615 = 8'h67 == req_index ? dirty_103 : _GEN_614; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_616 = 8'h68 == req_index ? dirty_104 : _GEN_615; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_617 = 8'h69 == req_index ? dirty_105 : _GEN_616; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_618 = 8'h6a == req_index ? dirty_106 : _GEN_617; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_619 = 8'h6b == req_index ? dirty_107 : _GEN_618; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_620 = 8'h6c == req_index ? dirty_108 : _GEN_619; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_621 = 8'h6d == req_index ? dirty_109 : _GEN_620; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_622 = 8'h6e == req_index ? dirty_110 : _GEN_621; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_623 = 8'h6f == req_index ? dirty_111 : _GEN_622; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_624 = 8'h70 == req_index ? dirty_112 : _GEN_623; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_625 = 8'h71 == req_index ? dirty_113 : _GEN_624; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_626 = 8'h72 == req_index ? dirty_114 : _GEN_625; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_627 = 8'h73 == req_index ? dirty_115 : _GEN_626; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_628 = 8'h74 == req_index ? dirty_116 : _GEN_627; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_629 = 8'h75 == req_index ? dirty_117 : _GEN_628; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_630 = 8'h76 == req_index ? dirty_118 : _GEN_629; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_631 = 8'h77 == req_index ? dirty_119 : _GEN_630; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_632 = 8'h78 == req_index ? dirty_120 : _GEN_631; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_633 = 8'h79 == req_index ? dirty_121 : _GEN_632; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_634 = 8'h7a == req_index ? dirty_122 : _GEN_633; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_635 = 8'h7b == req_index ? dirty_123 : _GEN_634; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_636 = 8'h7c == req_index ? dirty_124 : _GEN_635; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_637 = 8'h7d == req_index ? dirty_125 : _GEN_636; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_638 = 8'h7e == req_index ? dirty_126 : _GEN_637; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_639 = 8'h7f == req_index ? dirty_127 : _GEN_638; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_640 = 8'h80 == req_index ? dirty_128 : _GEN_639; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_641 = 8'h81 == req_index ? dirty_129 : _GEN_640; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_642 = 8'h82 == req_index ? dirty_130 : _GEN_641; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_643 = 8'h83 == req_index ? dirty_131 : _GEN_642; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_644 = 8'h84 == req_index ? dirty_132 : _GEN_643; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_645 = 8'h85 == req_index ? dirty_133 : _GEN_644; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_646 = 8'h86 == req_index ? dirty_134 : _GEN_645; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_647 = 8'h87 == req_index ? dirty_135 : _GEN_646; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_648 = 8'h88 == req_index ? dirty_136 : _GEN_647; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_649 = 8'h89 == req_index ? dirty_137 : _GEN_648; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_650 = 8'h8a == req_index ? dirty_138 : _GEN_649; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_651 = 8'h8b == req_index ? dirty_139 : _GEN_650; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_652 = 8'h8c == req_index ? dirty_140 : _GEN_651; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_653 = 8'h8d == req_index ? dirty_141 : _GEN_652; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_654 = 8'h8e == req_index ? dirty_142 : _GEN_653; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_655 = 8'h8f == req_index ? dirty_143 : _GEN_654; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_656 = 8'h90 == req_index ? dirty_144 : _GEN_655; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_657 = 8'h91 == req_index ? dirty_145 : _GEN_656; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_658 = 8'h92 == req_index ? dirty_146 : _GEN_657; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_659 = 8'h93 == req_index ? dirty_147 : _GEN_658; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_660 = 8'h94 == req_index ? dirty_148 : _GEN_659; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_661 = 8'h95 == req_index ? dirty_149 : _GEN_660; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_662 = 8'h96 == req_index ? dirty_150 : _GEN_661; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_663 = 8'h97 == req_index ? dirty_151 : _GEN_662; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_664 = 8'h98 == req_index ? dirty_152 : _GEN_663; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_665 = 8'h99 == req_index ? dirty_153 : _GEN_664; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_666 = 8'h9a == req_index ? dirty_154 : _GEN_665; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_667 = 8'h9b == req_index ? dirty_155 : _GEN_666; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_668 = 8'h9c == req_index ? dirty_156 : _GEN_667; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_669 = 8'h9d == req_index ? dirty_157 : _GEN_668; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_670 = 8'h9e == req_index ? dirty_158 : _GEN_669; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_671 = 8'h9f == req_index ? dirty_159 : _GEN_670; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_672 = 8'ha0 == req_index ? dirty_160 : _GEN_671; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_673 = 8'ha1 == req_index ? dirty_161 : _GEN_672; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_674 = 8'ha2 == req_index ? dirty_162 : _GEN_673; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_675 = 8'ha3 == req_index ? dirty_163 : _GEN_674; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_676 = 8'ha4 == req_index ? dirty_164 : _GEN_675; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_677 = 8'ha5 == req_index ? dirty_165 : _GEN_676; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_678 = 8'ha6 == req_index ? dirty_166 : _GEN_677; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_679 = 8'ha7 == req_index ? dirty_167 : _GEN_678; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_680 = 8'ha8 == req_index ? dirty_168 : _GEN_679; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_681 = 8'ha9 == req_index ? dirty_169 : _GEN_680; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_682 = 8'haa == req_index ? dirty_170 : _GEN_681; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_683 = 8'hab == req_index ? dirty_171 : _GEN_682; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_684 = 8'hac == req_index ? dirty_172 : _GEN_683; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_685 = 8'had == req_index ? dirty_173 : _GEN_684; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_686 = 8'hae == req_index ? dirty_174 : _GEN_685; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_687 = 8'haf == req_index ? dirty_175 : _GEN_686; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_688 = 8'hb0 == req_index ? dirty_176 : _GEN_687; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_689 = 8'hb1 == req_index ? dirty_177 : _GEN_688; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_690 = 8'hb2 == req_index ? dirty_178 : _GEN_689; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_691 = 8'hb3 == req_index ? dirty_179 : _GEN_690; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_692 = 8'hb4 == req_index ? dirty_180 : _GEN_691; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_693 = 8'hb5 == req_index ? dirty_181 : _GEN_692; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_694 = 8'hb6 == req_index ? dirty_182 : _GEN_693; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_695 = 8'hb7 == req_index ? dirty_183 : _GEN_694; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_696 = 8'hb8 == req_index ? dirty_184 : _GEN_695; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_697 = 8'hb9 == req_index ? dirty_185 : _GEN_696; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_698 = 8'hba == req_index ? dirty_186 : _GEN_697; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_699 = 8'hbb == req_index ? dirty_187 : _GEN_698; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_700 = 8'hbc == req_index ? dirty_188 : _GEN_699; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_701 = 8'hbd == req_index ? dirty_189 : _GEN_700; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_702 = 8'hbe == req_index ? dirty_190 : _GEN_701; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_703 = 8'hbf == req_index ? dirty_191 : _GEN_702; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_704 = 8'hc0 == req_index ? dirty_192 : _GEN_703; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_705 = 8'hc1 == req_index ? dirty_193 : _GEN_704; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_706 = 8'hc2 == req_index ? dirty_194 : _GEN_705; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_707 = 8'hc3 == req_index ? dirty_195 : _GEN_706; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_708 = 8'hc4 == req_index ? dirty_196 : _GEN_707; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_709 = 8'hc5 == req_index ? dirty_197 : _GEN_708; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_710 = 8'hc6 == req_index ? dirty_198 : _GEN_709; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_711 = 8'hc7 == req_index ? dirty_199 : _GEN_710; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_712 = 8'hc8 == req_index ? dirty_200 : _GEN_711; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_713 = 8'hc9 == req_index ? dirty_201 : _GEN_712; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_714 = 8'hca == req_index ? dirty_202 : _GEN_713; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_715 = 8'hcb == req_index ? dirty_203 : _GEN_714; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_716 = 8'hcc == req_index ? dirty_204 : _GEN_715; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_717 = 8'hcd == req_index ? dirty_205 : _GEN_716; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_718 = 8'hce == req_index ? dirty_206 : _GEN_717; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_719 = 8'hcf == req_index ? dirty_207 : _GEN_718; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_720 = 8'hd0 == req_index ? dirty_208 : _GEN_719; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_721 = 8'hd1 == req_index ? dirty_209 : _GEN_720; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_722 = 8'hd2 == req_index ? dirty_210 : _GEN_721; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_723 = 8'hd3 == req_index ? dirty_211 : _GEN_722; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_724 = 8'hd4 == req_index ? dirty_212 : _GEN_723; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_725 = 8'hd5 == req_index ? dirty_213 : _GEN_724; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_726 = 8'hd6 == req_index ? dirty_214 : _GEN_725; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_727 = 8'hd7 == req_index ? dirty_215 : _GEN_726; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_728 = 8'hd8 == req_index ? dirty_216 : _GEN_727; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_729 = 8'hd9 == req_index ? dirty_217 : _GEN_728; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_730 = 8'hda == req_index ? dirty_218 : _GEN_729; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_731 = 8'hdb == req_index ? dirty_219 : _GEN_730; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_732 = 8'hdc == req_index ? dirty_220 : _GEN_731; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_733 = 8'hdd == req_index ? dirty_221 : _GEN_732; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_734 = 8'hde == req_index ? dirty_222 : _GEN_733; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_735 = 8'hdf == req_index ? dirty_223 : _GEN_734; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_736 = 8'he0 == req_index ? dirty_224 : _GEN_735; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_737 = 8'he1 == req_index ? dirty_225 : _GEN_736; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_738 = 8'he2 == req_index ? dirty_226 : _GEN_737; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_739 = 8'he3 == req_index ? dirty_227 : _GEN_738; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_740 = 8'he4 == req_index ? dirty_228 : _GEN_739; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_741 = 8'he5 == req_index ? dirty_229 : _GEN_740; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_742 = 8'he6 == req_index ? dirty_230 : _GEN_741; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_743 = 8'he7 == req_index ? dirty_231 : _GEN_742; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_744 = 8'he8 == req_index ? dirty_232 : _GEN_743; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_745 = 8'he9 == req_index ? dirty_233 : _GEN_744; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_746 = 8'hea == req_index ? dirty_234 : _GEN_745; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_747 = 8'heb == req_index ? dirty_235 : _GEN_746; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_748 = 8'hec == req_index ? dirty_236 : _GEN_747; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_749 = 8'hed == req_index ? dirty_237 : _GEN_748; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_750 = 8'hee == req_index ? dirty_238 : _GEN_749; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_751 = 8'hef == req_index ? dirty_239 : _GEN_750; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_752 = 8'hf0 == req_index ? dirty_240 : _GEN_751; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_753 = 8'hf1 == req_index ? dirty_241 : _GEN_752; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_754 = 8'hf2 == req_index ? dirty_242 : _GEN_753; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_755 = 8'hf3 == req_index ? dirty_243 : _GEN_754; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_756 = 8'hf4 == req_index ? dirty_244 : _GEN_755; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_757 = 8'hf5 == req_index ? dirty_245 : _GEN_756; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_758 = 8'hf6 == req_index ? dirty_246 : _GEN_757; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_759 = 8'hf7 == req_index ? dirty_247 : _GEN_758; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_760 = 8'hf8 == req_index ? dirty_248 : _GEN_759; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_761 = 8'hf9 == req_index ? dirty_249 : _GEN_760; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_762 = 8'hfa == req_index ? dirty_250 : _GEN_761; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_763 = 8'hfb == req_index ? dirty_251 : _GEN_762; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_764 = 8'hfc == req_index ? dirty_252 : _GEN_763; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_765 = 8'hfd == req_index ? dirty_253 : _GEN_764; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_766 = 8'hfe == req_index ? dirty_254 : _GEN_765; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_767 = 8'hff == req_index ? dirty_255 : _GEN_766; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  cache_dirty = _GEN_767 & _cache_hit_T_2; // @[Dcache.scala 35:38]
  reg  data_ready; // @[Dcache.scala 46:28]
  wire [127:0] cache_data_out = req_Q; // @[Dcache.scala 37:28 Dcache.scala 227:18]
  wire [63:0] valid_rdata = req_offset[3] ? cache_data_out[127:64] : cache_data_out[63:0]; // @[Dcache.scala 48:24]
  wire [7:0] _valid_strb_T_1 = 8'h1 == io_dmem_data_strb ? 8'hff : 8'h0; // @[Mux.scala 80:57]
  wire [15:0] _valid_strb_T_3 = 8'h2 == io_dmem_data_strb ? 16'hff00 : {{8'd0}, _valid_strb_T_1}; // @[Mux.scala 80:57]
  wire [23:0] _valid_strb_T_5 = 8'h4 == io_dmem_data_strb ? 24'hff0000 : {{8'd0}, _valid_strb_T_3}; // @[Mux.scala 80:57]
  wire [31:0] _valid_strb_T_7 = 8'h8 == io_dmem_data_strb ? 32'hff000000 : {{8'd0}, _valid_strb_T_5}; // @[Mux.scala 80:57]
  wire [39:0] _valid_strb_T_9 = 8'h10 == io_dmem_data_strb ? 40'hff00000000 : {{8'd0}, _valid_strb_T_7}; // @[Mux.scala 80:57]
  wire [47:0] _valid_strb_T_11 = 8'h20 == io_dmem_data_strb ? 48'hff0000000000 : {{8'd0}, _valid_strb_T_9}; // @[Mux.scala 80:57]
  wire [55:0] _valid_strb_T_13 = 8'h40 == io_dmem_data_strb ? 56'hff000000000000 : {{8'd0}, _valid_strb_T_11}; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_15 = 8'h80 == io_dmem_data_strb ? 64'hff00000000000000 : {{8'd0}, _valid_strb_T_13}; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_17 = 8'h3 == io_dmem_data_strb ? 64'hffff : _valid_strb_T_15; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_19 = 8'hc == io_dmem_data_strb ? 64'hffff0000 : _valid_strb_T_17; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_21 = 8'h30 == io_dmem_data_strb ? 64'hffff00000000 : _valid_strb_T_19; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_23 = 8'hc0 == io_dmem_data_strb ? 64'hffff000000000000 : _valid_strb_T_21; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_25 = 8'hf == io_dmem_data_strb ? 64'hffffffff : _valid_strb_T_23; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_27 = 8'hf0 == io_dmem_data_strb ? 64'hffffffff00000000 : _valid_strb_T_25; // @[Mux.scala 80:57]
  wire [63:0] valid_strb = 8'hff == io_dmem_data_strb ? 64'hffffffffffffffff : _valid_strb_T_27; // @[Mux.scala 80:57]
  wire [63:0] valid_data = req_offset[3] ? io_out_data_read[127:64] : io_out_data_read[63:0]; // @[Dcache.scala 67:24]
  wire [55:0] valid_wdata_hi = valid_data[63:8]; // @[Dcache.scala 70:47]
  wire [7:0] valid_wdata_lo = io_dmem_data_write[7:0]; // @[Dcache.scala 70:69]
  wire [63:0] _valid_wdata_T_1 = {valid_wdata_hi,valid_wdata_lo}; // @[Cat.scala 30:58]
  wire [47:0] valid_wdata_hi_hi = valid_data[63:16]; // @[Dcache.scala 71:47]
  wire [7:0] valid_wdata_hi_lo = io_dmem_data_write[15:8]; // @[Dcache.scala 71:69]
  wire [7:0] valid_wdata_lo_1 = valid_data[7:0]; // @[Dcache.scala 71:88]
  wire [63:0] _valid_wdata_T_2 = {valid_wdata_hi_hi,valid_wdata_hi_lo,valid_wdata_lo_1}; // @[Cat.scala 30:58]
  wire [39:0] valid_wdata_hi_hi_1 = valid_data[63:24]; // @[Dcache.scala 72:47]
  wire [7:0] valid_wdata_hi_lo_1 = io_dmem_data_write[23:16]; // @[Dcache.scala 72:69]
  wire [15:0] valid_wdata_lo_2 = valid_data[15:0]; // @[Dcache.scala 72:88]
  wire [63:0] _valid_wdata_T_3 = {valid_wdata_hi_hi_1,valid_wdata_hi_lo_1,valid_wdata_lo_2}; // @[Cat.scala 30:58]
  wire [31:0] valid_wdata_hi_hi_2 = valid_data[63:32]; // @[Dcache.scala 73:47]
  wire [7:0] valid_wdata_hi_lo_2 = io_dmem_data_write[31:24]; // @[Dcache.scala 73:69]
  wire [23:0] valid_wdata_lo_3 = valid_data[23:0]; // @[Dcache.scala 73:88]
  wire [63:0] _valid_wdata_T_4 = {valid_wdata_hi_hi_2,valid_wdata_hi_lo_2,valid_wdata_lo_3}; // @[Cat.scala 30:58]
  wire [23:0] valid_wdata_hi_hi_3 = valid_data[63:40]; // @[Dcache.scala 74:47]
  wire [7:0] valid_wdata_hi_lo_3 = io_dmem_data_write[39:32]; // @[Dcache.scala 74:69]
  wire [31:0] valid_wdata_lo_4 = valid_data[31:0]; // @[Dcache.scala 74:88]
  wire [63:0] _valid_wdata_T_5 = {valid_wdata_hi_hi_3,valid_wdata_hi_lo_3,valid_wdata_lo_4}; // @[Cat.scala 30:58]
  wire [15:0] valid_wdata_hi_hi_4 = valid_data[63:48]; // @[Dcache.scala 75:47]
  wire [7:0] valid_wdata_hi_lo_4 = io_dmem_data_write[47:40]; // @[Dcache.scala 75:69]
  wire [39:0] valid_wdata_lo_5 = valid_data[39:0]; // @[Dcache.scala 75:88]
  wire [63:0] _valid_wdata_T_6 = {valid_wdata_hi_hi_4,valid_wdata_hi_lo_4,valid_wdata_lo_5}; // @[Cat.scala 30:58]
  wire [7:0] valid_wdata_hi_hi_5 = valid_data[63:56]; // @[Dcache.scala 76:47]
  wire [7:0] valid_wdata_hi_lo_5 = io_dmem_data_write[55:48]; // @[Dcache.scala 76:69]
  wire [47:0] valid_wdata_lo_6 = valid_data[47:0]; // @[Dcache.scala 76:88]
  wire [63:0] _valid_wdata_T_7 = {valid_wdata_hi_hi_5,valid_wdata_hi_lo_5,valid_wdata_lo_6}; // @[Cat.scala 30:58]
  wire [7:0] valid_wdata_hi_7 = io_dmem_data_write[63:56]; // @[Dcache.scala 77:50]
  wire [55:0] valid_wdata_lo_7 = valid_data[55:0]; // @[Dcache.scala 77:69]
  wire [63:0] _valid_wdata_T_8 = {valid_wdata_hi_7,valid_wdata_lo_7}; // @[Cat.scala 30:58]
  wire [63:0] _valid_wdata_T_10 = 3'h1 == req_offset[2:0] ? _valid_wdata_T_2 : _valid_wdata_T_1; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_12 = 3'h2 == req_offset[2:0] ? _valid_wdata_T_3 : _valid_wdata_T_10; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_14 = 3'h3 == req_offset[2:0] ? _valid_wdata_T_4 : _valid_wdata_T_12; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_16 = 3'h4 == req_offset[2:0] ? _valid_wdata_T_5 : _valid_wdata_T_14; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_18 = 3'h5 == req_offset[2:0] ? _valid_wdata_T_6 : _valid_wdata_T_16; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_20 = 3'h6 == req_offset[2:0] ? _valid_wdata_T_7 : _valid_wdata_T_18; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_22 = 3'h7 == req_offset[2:0] ? _valid_wdata_T_8 : _valid_wdata_T_20; // @[Mux.scala 80:57]
  wire [15:0] valid_wdata_lo_8 = io_dmem_data_write[15:0]; // @[Dcache.scala 80:68]
  wire [63:0] _valid_wdata_T_24 = {valid_wdata_hi_hi,valid_wdata_lo_8}; // @[Cat.scala 30:58]
  wire [15:0] valid_wdata_hi_lo_6 = io_dmem_data_write[31:16]; // @[Dcache.scala 81:68]
  wire [63:0] _valid_wdata_T_25 = {valid_wdata_hi_hi_2,valid_wdata_hi_lo_6,valid_wdata_lo_2}; // @[Cat.scala 30:58]
  wire [15:0] valid_wdata_hi_lo_7 = io_dmem_data_write[47:32]; // @[Dcache.scala 82:68]
  wire [63:0] _valid_wdata_T_26 = {valid_wdata_hi_hi_4,valid_wdata_hi_lo_7,valid_wdata_lo_4}; // @[Cat.scala 30:58]
  wire [15:0] valid_wdata_hi_11 = io_dmem_data_write[63:48]; // @[Dcache.scala 83:49]
  wire [63:0] _valid_wdata_T_27 = {valid_wdata_hi_11,valid_wdata_lo_6}; // @[Cat.scala 30:58]
  wire [63:0] _valid_wdata_T_29 = 2'h1 == req_offset[2:1] ? _valid_wdata_T_25 : _valid_wdata_T_24; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_31 = 2'h2 == req_offset[2:1] ? _valid_wdata_T_26 : _valid_wdata_T_29; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_33 = 2'h3 == req_offset[2:1] ? _valid_wdata_T_27 : _valid_wdata_T_31; // @[Mux.scala 80:57]
  wire [31:0] valid_wdata_lo_12 = io_dmem_data_write[31:0]; // @[Dcache.scala 86:67]
  wire [63:0] _valid_wdata_T_35 = {valid_wdata_hi_hi_2,valid_wdata_lo_12}; // @[Cat.scala 30:58]
  wire [31:0] valid_wdata_hi_13 = io_dmem_data_write[63:32]; // @[Dcache.scala 87:48]
  wire [63:0] _valid_wdata_T_36 = {valid_wdata_hi_13,valid_wdata_lo_4}; // @[Cat.scala 30:58]
  wire [63:0] _valid_wdata_T_38 = req_offset[2] ? _valid_wdata_T_36 : _valid_wdata_T_35; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_40 = 2'h1 == io_dmem_data_size ? _valid_wdata_T_33 : _valid_wdata_T_22; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_42 = 2'h2 == io_dmem_data_size ? _valid_wdata_T_38 : _valid_wdata_T_40; // @[Mux.scala 80:57]
  wire [63:0] valid_wdata = 2'h3 == io_dmem_data_size ? io_dmem_data_write : _valid_wdata_T_42; // @[Mux.scala 80:57]
  wire [7:0] data_read_lo = valid_rdata[7:0]; // @[Dcache.scala 94:53]
  wire [8:0] _data_read_T_1 = {1'h0,data_read_lo}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_1 = valid_rdata[15:8]; // @[Dcache.scala 95:53]
  wire [8:0] _data_read_T_2 = {1'h0,data_read_lo_1}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_2 = valid_rdata[23:16]; // @[Dcache.scala 96:53]
  wire [8:0] _data_read_T_3 = {1'h0,data_read_lo_2}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_3 = valid_rdata[31:24]; // @[Dcache.scala 97:53]
  wire [8:0] _data_read_T_4 = {1'h0,data_read_lo_3}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_4 = valid_rdata[39:32]; // @[Dcache.scala 98:53]
  wire [8:0] _data_read_T_5 = {1'h0,data_read_lo_4}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_5 = valid_rdata[47:40]; // @[Dcache.scala 99:53]
  wire [8:0] _data_read_T_6 = {1'h0,data_read_lo_5}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_6 = valid_rdata[55:48]; // @[Dcache.scala 100:53]
  wire [8:0] _data_read_T_7 = {1'h0,data_read_lo_6}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_7 = valid_rdata[63:56]; // @[Dcache.scala 101:53]
  wire [8:0] _data_read_T_8 = {1'h0,data_read_lo_7}; // @[Cat.scala 30:58]
  wire [8:0] _data_read_T_10 = 3'h1 == req_offset[2:0] ? _data_read_T_2 : _data_read_T_1; // @[Mux.scala 80:57]
  wire [8:0] _data_read_T_12 = 3'h2 == req_offset[2:0] ? _data_read_T_3 : _data_read_T_10; // @[Mux.scala 80:57]
  wire [8:0] _data_read_T_14 = 3'h3 == req_offset[2:0] ? _data_read_T_4 : _data_read_T_12; // @[Mux.scala 80:57]
  wire [8:0] _data_read_T_16 = 3'h4 == req_offset[2:0] ? _data_read_T_5 : _data_read_T_14; // @[Mux.scala 80:57]
  wire [8:0] _data_read_T_18 = 3'h5 == req_offset[2:0] ? _data_read_T_6 : _data_read_T_16; // @[Mux.scala 80:57]
  wire [8:0] _data_read_T_20 = 3'h6 == req_offset[2:0] ? _data_read_T_7 : _data_read_T_18; // @[Mux.scala 80:57]
  wire [8:0] _data_read_T_22 = 3'h7 == req_offset[2:0] ? _data_read_T_8 : _data_read_T_20; // @[Mux.scala 80:57]
  wire [15:0] data_read_lo_8 = valid_rdata[15:0]; // @[Dcache.scala 104:52]
  wire [16:0] _data_read_T_24 = {1'h0,data_read_lo_8}; // @[Cat.scala 30:58]
  wire [15:0] data_read_lo_9 = valid_rdata[31:16]; // @[Dcache.scala 105:52]
  wire [16:0] _data_read_T_25 = {1'h0,data_read_lo_9}; // @[Cat.scala 30:58]
  wire [15:0] data_read_lo_10 = valid_rdata[47:32]; // @[Dcache.scala 106:52]
  wire [16:0] _data_read_T_26 = {1'h0,data_read_lo_10}; // @[Cat.scala 30:58]
  wire [15:0] data_read_lo_11 = valid_rdata[63:48]; // @[Dcache.scala 107:52]
  wire [16:0] _data_read_T_27 = {1'h0,data_read_lo_11}; // @[Cat.scala 30:58]
  wire [16:0] _data_read_T_29 = 2'h1 == req_offset[2:1] ? _data_read_T_25 : _data_read_T_24; // @[Mux.scala 80:57]
  wire [16:0] _data_read_T_31 = 2'h2 == req_offset[2:1] ? _data_read_T_26 : _data_read_T_29; // @[Mux.scala 80:57]
  wire [16:0] _data_read_T_33 = 2'h3 == req_offset[2:1] ? _data_read_T_27 : _data_read_T_31; // @[Mux.scala 80:57]
  wire [31:0] data_read_lo_12 = valid_rdata[31:0]; // @[Dcache.scala 110:51]
  wire [32:0] _data_read_T_35 = {1'h0,data_read_lo_12}; // @[Cat.scala 30:58]
  wire [31:0] data_read_lo_13 = valid_rdata[63:32]; // @[Dcache.scala 111:51]
  wire [32:0] _data_read_T_36 = {1'h0,data_read_lo_13}; // @[Cat.scala 30:58]
  wire [32:0] _data_read_T_38 = req_offset[2] ? _data_read_T_36 : _data_read_T_35; // @[Mux.scala 80:57]
  wire [16:0] _data_read_T_40 = 2'h1 == io_dmem_data_size ? _data_read_T_33 : {{8'd0}, _data_read_T_22}; // @[Mux.scala 80:57]
  wire [32:0] _data_read_T_42 = 2'h2 == io_dmem_data_size ? _data_read_T_38 : {{16'd0}, _data_read_T_40}; // @[Mux.scala 80:57]
  reg  cache_fill; // @[Dcache.scala 116:28]
  reg  cache_wen; // @[Dcache.scala 117:28]
  reg [127:0] cache_wdata; // @[Dcache.scala 118:28]
  reg [127:0] cache_strb; // @[Dcache.scala 119:28]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _GEN_769 = 8'h0 == req_index | valid_0; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_770 = 8'h1 == req_index | valid_1; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_771 = 8'h2 == req_index | valid_2; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_772 = 8'h3 == req_index | valid_3; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_773 = 8'h4 == req_index | valid_4; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_774 = 8'h5 == req_index | valid_5; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_775 = 8'h6 == req_index | valid_6; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_776 = 8'h7 == req_index | valid_7; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_777 = 8'h8 == req_index | valid_8; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_778 = 8'h9 == req_index | valid_9; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_779 = 8'ha == req_index | valid_10; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_780 = 8'hb == req_index | valid_11; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_781 = 8'hc == req_index | valid_12; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_782 = 8'hd == req_index | valid_13; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_783 = 8'he == req_index | valid_14; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_784 = 8'hf == req_index | valid_15; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_785 = 8'h10 == req_index | valid_16; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_786 = 8'h11 == req_index | valid_17; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_787 = 8'h12 == req_index | valid_18; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_788 = 8'h13 == req_index | valid_19; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_789 = 8'h14 == req_index | valid_20; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_790 = 8'h15 == req_index | valid_21; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_791 = 8'h16 == req_index | valid_22; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_792 = 8'h17 == req_index | valid_23; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_793 = 8'h18 == req_index | valid_24; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_794 = 8'h19 == req_index | valid_25; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_795 = 8'h1a == req_index | valid_26; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_796 = 8'h1b == req_index | valid_27; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_797 = 8'h1c == req_index | valid_28; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_798 = 8'h1d == req_index | valid_29; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_799 = 8'h1e == req_index | valid_30; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_800 = 8'h1f == req_index | valid_31; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_801 = 8'h20 == req_index | valid_32; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_802 = 8'h21 == req_index | valid_33; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_803 = 8'h22 == req_index | valid_34; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_804 = 8'h23 == req_index | valid_35; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_805 = 8'h24 == req_index | valid_36; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_806 = 8'h25 == req_index | valid_37; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_807 = 8'h26 == req_index | valid_38; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_808 = 8'h27 == req_index | valid_39; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_809 = 8'h28 == req_index | valid_40; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_810 = 8'h29 == req_index | valid_41; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_811 = 8'h2a == req_index | valid_42; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_812 = 8'h2b == req_index | valid_43; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_813 = 8'h2c == req_index | valid_44; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_814 = 8'h2d == req_index | valid_45; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_815 = 8'h2e == req_index | valid_46; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_816 = 8'h2f == req_index | valid_47; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_817 = 8'h30 == req_index | valid_48; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_818 = 8'h31 == req_index | valid_49; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_819 = 8'h32 == req_index | valid_50; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_820 = 8'h33 == req_index | valid_51; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_821 = 8'h34 == req_index | valid_52; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_822 = 8'h35 == req_index | valid_53; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_823 = 8'h36 == req_index | valid_54; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_824 = 8'h37 == req_index | valid_55; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_825 = 8'h38 == req_index | valid_56; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_826 = 8'h39 == req_index | valid_57; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_827 = 8'h3a == req_index | valid_58; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_828 = 8'h3b == req_index | valid_59; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_829 = 8'h3c == req_index | valid_60; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_830 = 8'h3d == req_index | valid_61; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_831 = 8'h3e == req_index | valid_62; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_832 = 8'h3f == req_index | valid_63; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_833 = 8'h40 == req_index | valid_64; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_834 = 8'h41 == req_index | valid_65; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_835 = 8'h42 == req_index | valid_66; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_836 = 8'h43 == req_index | valid_67; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_837 = 8'h44 == req_index | valid_68; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_838 = 8'h45 == req_index | valid_69; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_839 = 8'h46 == req_index | valid_70; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_840 = 8'h47 == req_index | valid_71; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_841 = 8'h48 == req_index | valid_72; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_842 = 8'h49 == req_index | valid_73; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_843 = 8'h4a == req_index | valid_74; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_844 = 8'h4b == req_index | valid_75; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_845 = 8'h4c == req_index | valid_76; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_846 = 8'h4d == req_index | valid_77; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_847 = 8'h4e == req_index | valid_78; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_848 = 8'h4f == req_index | valid_79; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_849 = 8'h50 == req_index | valid_80; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_850 = 8'h51 == req_index | valid_81; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_851 = 8'h52 == req_index | valid_82; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_852 = 8'h53 == req_index | valid_83; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_853 = 8'h54 == req_index | valid_84; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_854 = 8'h55 == req_index | valid_85; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_855 = 8'h56 == req_index | valid_86; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_856 = 8'h57 == req_index | valid_87; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_857 = 8'h58 == req_index | valid_88; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_858 = 8'h59 == req_index | valid_89; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_859 = 8'h5a == req_index | valid_90; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_860 = 8'h5b == req_index | valid_91; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_861 = 8'h5c == req_index | valid_92; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_862 = 8'h5d == req_index | valid_93; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_863 = 8'h5e == req_index | valid_94; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_864 = 8'h5f == req_index | valid_95; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_865 = 8'h60 == req_index | valid_96; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_866 = 8'h61 == req_index | valid_97; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_867 = 8'h62 == req_index | valid_98; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_868 = 8'h63 == req_index | valid_99; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_869 = 8'h64 == req_index | valid_100; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_870 = 8'h65 == req_index | valid_101; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_871 = 8'h66 == req_index | valid_102; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_872 = 8'h67 == req_index | valid_103; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_873 = 8'h68 == req_index | valid_104; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_874 = 8'h69 == req_index | valid_105; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_875 = 8'h6a == req_index | valid_106; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_876 = 8'h6b == req_index | valid_107; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_877 = 8'h6c == req_index | valid_108; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_878 = 8'h6d == req_index | valid_109; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_879 = 8'h6e == req_index | valid_110; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_880 = 8'h6f == req_index | valid_111; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_881 = 8'h70 == req_index | valid_112; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_882 = 8'h71 == req_index | valid_113; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_883 = 8'h72 == req_index | valid_114; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_884 = 8'h73 == req_index | valid_115; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_885 = 8'h74 == req_index | valid_116; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_886 = 8'h75 == req_index | valid_117; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_887 = 8'h76 == req_index | valid_118; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_888 = 8'h77 == req_index | valid_119; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_889 = 8'h78 == req_index | valid_120; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_890 = 8'h79 == req_index | valid_121; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_891 = 8'h7a == req_index | valid_122; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_892 = 8'h7b == req_index | valid_123; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_893 = 8'h7c == req_index | valid_124; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_894 = 8'h7d == req_index | valid_125; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_895 = 8'h7e == req_index | valid_126; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_896 = 8'h7f == req_index | valid_127; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_897 = 8'h80 == req_index | valid_128; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_898 = 8'h81 == req_index | valid_129; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_899 = 8'h82 == req_index | valid_130; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_900 = 8'h83 == req_index | valid_131; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_901 = 8'h84 == req_index | valid_132; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_902 = 8'h85 == req_index | valid_133; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_903 = 8'h86 == req_index | valid_134; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_904 = 8'h87 == req_index | valid_135; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_905 = 8'h88 == req_index | valid_136; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_906 = 8'h89 == req_index | valid_137; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_907 = 8'h8a == req_index | valid_138; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_908 = 8'h8b == req_index | valid_139; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_909 = 8'h8c == req_index | valid_140; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_910 = 8'h8d == req_index | valid_141; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_911 = 8'h8e == req_index | valid_142; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_912 = 8'h8f == req_index | valid_143; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_913 = 8'h90 == req_index | valid_144; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_914 = 8'h91 == req_index | valid_145; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_915 = 8'h92 == req_index | valid_146; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_916 = 8'h93 == req_index | valid_147; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_917 = 8'h94 == req_index | valid_148; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_918 = 8'h95 == req_index | valid_149; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_919 = 8'h96 == req_index | valid_150; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_920 = 8'h97 == req_index | valid_151; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_921 = 8'h98 == req_index | valid_152; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_922 = 8'h99 == req_index | valid_153; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_923 = 8'h9a == req_index | valid_154; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_924 = 8'h9b == req_index | valid_155; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_925 = 8'h9c == req_index | valid_156; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_926 = 8'h9d == req_index | valid_157; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_927 = 8'h9e == req_index | valid_158; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_928 = 8'h9f == req_index | valid_159; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_929 = 8'ha0 == req_index | valid_160; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_930 = 8'ha1 == req_index | valid_161; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_931 = 8'ha2 == req_index | valid_162; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_932 = 8'ha3 == req_index | valid_163; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_933 = 8'ha4 == req_index | valid_164; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_934 = 8'ha5 == req_index | valid_165; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_935 = 8'ha6 == req_index | valid_166; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_936 = 8'ha7 == req_index | valid_167; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_937 = 8'ha8 == req_index | valid_168; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_938 = 8'ha9 == req_index | valid_169; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_939 = 8'haa == req_index | valid_170; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_940 = 8'hab == req_index | valid_171; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_941 = 8'hac == req_index | valid_172; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_942 = 8'had == req_index | valid_173; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_943 = 8'hae == req_index | valid_174; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_944 = 8'haf == req_index | valid_175; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_945 = 8'hb0 == req_index | valid_176; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_946 = 8'hb1 == req_index | valid_177; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_947 = 8'hb2 == req_index | valid_178; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_948 = 8'hb3 == req_index | valid_179; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_949 = 8'hb4 == req_index | valid_180; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_950 = 8'hb5 == req_index | valid_181; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_951 = 8'hb6 == req_index | valid_182; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_952 = 8'hb7 == req_index | valid_183; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_953 = 8'hb8 == req_index | valid_184; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_954 = 8'hb9 == req_index | valid_185; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_955 = 8'hba == req_index | valid_186; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_956 = 8'hbb == req_index | valid_187; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_957 = 8'hbc == req_index | valid_188; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_958 = 8'hbd == req_index | valid_189; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_959 = 8'hbe == req_index | valid_190; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_960 = 8'hbf == req_index | valid_191; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_961 = 8'hc0 == req_index | valid_192; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_962 = 8'hc1 == req_index | valid_193; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_963 = 8'hc2 == req_index | valid_194; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_964 = 8'hc3 == req_index | valid_195; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_965 = 8'hc4 == req_index | valid_196; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_966 = 8'hc5 == req_index | valid_197; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_967 = 8'hc6 == req_index | valid_198; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_968 = 8'hc7 == req_index | valid_199; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_969 = 8'hc8 == req_index | valid_200; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_970 = 8'hc9 == req_index | valid_201; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_971 = 8'hca == req_index | valid_202; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_972 = 8'hcb == req_index | valid_203; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_973 = 8'hcc == req_index | valid_204; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_974 = 8'hcd == req_index | valid_205; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_975 = 8'hce == req_index | valid_206; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_976 = 8'hcf == req_index | valid_207; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_977 = 8'hd0 == req_index | valid_208; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_978 = 8'hd1 == req_index | valid_209; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_979 = 8'hd2 == req_index | valid_210; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_980 = 8'hd3 == req_index | valid_211; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_981 = 8'hd4 == req_index | valid_212; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_982 = 8'hd5 == req_index | valid_213; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_983 = 8'hd6 == req_index | valid_214; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_984 = 8'hd7 == req_index | valid_215; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_985 = 8'hd8 == req_index | valid_216; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_986 = 8'hd9 == req_index | valid_217; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_987 = 8'hda == req_index | valid_218; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_988 = 8'hdb == req_index | valid_219; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_989 = 8'hdc == req_index | valid_220; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_990 = 8'hdd == req_index | valid_221; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_991 = 8'hde == req_index | valid_222; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_992 = 8'hdf == req_index | valid_223; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_993 = 8'he0 == req_index | valid_224; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_994 = 8'he1 == req_index | valid_225; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_995 = 8'he2 == req_index | valid_226; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_996 = 8'he3 == req_index | valid_227; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_997 = 8'he4 == req_index | valid_228; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_998 = 8'he5 == req_index | valid_229; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_999 = 8'he6 == req_index | valid_230; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1000 = 8'he7 == req_index | valid_231; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1001 = 8'he8 == req_index | valid_232; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1002 = 8'he9 == req_index | valid_233; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1003 = 8'hea == req_index | valid_234; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1004 = 8'heb == req_index | valid_235; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1005 = 8'hec == req_index | valid_236; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1006 = 8'hed == req_index | valid_237; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1007 = 8'hee == req_index | valid_238; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1008 = 8'hef == req_index | valid_239; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1009 = 8'hf0 == req_index | valid_240; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1010 = 8'hf1 == req_index | valid_241; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1011 = 8'hf2 == req_index | valid_242; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1012 = 8'hf3 == req_index | valid_243; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1013 = 8'hf4 == req_index | valid_244; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1014 = 8'hf5 == req_index | valid_245; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1015 = 8'hf6 == req_index | valid_246; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1016 = 8'hf7 == req_index | valid_247; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1017 = 8'hf8 == req_index | valid_248; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1018 = 8'hf9 == req_index | valid_249; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1019 = 8'hfa == req_index | valid_250; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1020 = 8'hfb == req_index | valid_251; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1021 = 8'hfc == req_index | valid_252; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1022 = 8'hfd == req_index | valid_253; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1023 = 8'hfe == req_index | valid_254; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire  _GEN_1024 = 8'hff == req_index | valid_255; // @[Dcache.scala 135:27 Dcache.scala 135:27 Dcache.scala 17:24]
  wire [19:0] _GEN_1025 = 8'h0 == req_index ? req_tag : tag_0; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1026 = 8'h1 == req_index ? req_tag : tag_1; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1027 = 8'h2 == req_index ? req_tag : tag_2; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1028 = 8'h3 == req_index ? req_tag : tag_3; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1029 = 8'h4 == req_index ? req_tag : tag_4; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1030 = 8'h5 == req_index ? req_tag : tag_5; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1031 = 8'h6 == req_index ? req_tag : tag_6; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1032 = 8'h7 == req_index ? req_tag : tag_7; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1033 = 8'h8 == req_index ? req_tag : tag_8; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1034 = 8'h9 == req_index ? req_tag : tag_9; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1035 = 8'ha == req_index ? req_tag : tag_10; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1036 = 8'hb == req_index ? req_tag : tag_11; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1037 = 8'hc == req_index ? req_tag : tag_12; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1038 = 8'hd == req_index ? req_tag : tag_13; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1039 = 8'he == req_index ? req_tag : tag_14; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1040 = 8'hf == req_index ? req_tag : tag_15; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1041 = 8'h10 == req_index ? req_tag : tag_16; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1042 = 8'h11 == req_index ? req_tag : tag_17; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1043 = 8'h12 == req_index ? req_tag : tag_18; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1044 = 8'h13 == req_index ? req_tag : tag_19; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1045 = 8'h14 == req_index ? req_tag : tag_20; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1046 = 8'h15 == req_index ? req_tag : tag_21; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1047 = 8'h16 == req_index ? req_tag : tag_22; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1048 = 8'h17 == req_index ? req_tag : tag_23; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1049 = 8'h18 == req_index ? req_tag : tag_24; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1050 = 8'h19 == req_index ? req_tag : tag_25; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1051 = 8'h1a == req_index ? req_tag : tag_26; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1052 = 8'h1b == req_index ? req_tag : tag_27; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1053 = 8'h1c == req_index ? req_tag : tag_28; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1054 = 8'h1d == req_index ? req_tag : tag_29; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1055 = 8'h1e == req_index ? req_tag : tag_30; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1056 = 8'h1f == req_index ? req_tag : tag_31; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1057 = 8'h20 == req_index ? req_tag : tag_32; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1058 = 8'h21 == req_index ? req_tag : tag_33; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1059 = 8'h22 == req_index ? req_tag : tag_34; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1060 = 8'h23 == req_index ? req_tag : tag_35; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1061 = 8'h24 == req_index ? req_tag : tag_36; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1062 = 8'h25 == req_index ? req_tag : tag_37; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1063 = 8'h26 == req_index ? req_tag : tag_38; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1064 = 8'h27 == req_index ? req_tag : tag_39; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1065 = 8'h28 == req_index ? req_tag : tag_40; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1066 = 8'h29 == req_index ? req_tag : tag_41; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1067 = 8'h2a == req_index ? req_tag : tag_42; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1068 = 8'h2b == req_index ? req_tag : tag_43; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1069 = 8'h2c == req_index ? req_tag : tag_44; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1070 = 8'h2d == req_index ? req_tag : tag_45; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1071 = 8'h2e == req_index ? req_tag : tag_46; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1072 = 8'h2f == req_index ? req_tag : tag_47; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1073 = 8'h30 == req_index ? req_tag : tag_48; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1074 = 8'h31 == req_index ? req_tag : tag_49; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1075 = 8'h32 == req_index ? req_tag : tag_50; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1076 = 8'h33 == req_index ? req_tag : tag_51; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1077 = 8'h34 == req_index ? req_tag : tag_52; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1078 = 8'h35 == req_index ? req_tag : tag_53; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1079 = 8'h36 == req_index ? req_tag : tag_54; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1080 = 8'h37 == req_index ? req_tag : tag_55; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1081 = 8'h38 == req_index ? req_tag : tag_56; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1082 = 8'h39 == req_index ? req_tag : tag_57; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1083 = 8'h3a == req_index ? req_tag : tag_58; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1084 = 8'h3b == req_index ? req_tag : tag_59; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1085 = 8'h3c == req_index ? req_tag : tag_60; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1086 = 8'h3d == req_index ? req_tag : tag_61; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1087 = 8'h3e == req_index ? req_tag : tag_62; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1088 = 8'h3f == req_index ? req_tag : tag_63; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1089 = 8'h40 == req_index ? req_tag : tag_64; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1090 = 8'h41 == req_index ? req_tag : tag_65; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1091 = 8'h42 == req_index ? req_tag : tag_66; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1092 = 8'h43 == req_index ? req_tag : tag_67; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1093 = 8'h44 == req_index ? req_tag : tag_68; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1094 = 8'h45 == req_index ? req_tag : tag_69; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1095 = 8'h46 == req_index ? req_tag : tag_70; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1096 = 8'h47 == req_index ? req_tag : tag_71; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1097 = 8'h48 == req_index ? req_tag : tag_72; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1098 = 8'h49 == req_index ? req_tag : tag_73; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1099 = 8'h4a == req_index ? req_tag : tag_74; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1100 = 8'h4b == req_index ? req_tag : tag_75; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1101 = 8'h4c == req_index ? req_tag : tag_76; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1102 = 8'h4d == req_index ? req_tag : tag_77; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1103 = 8'h4e == req_index ? req_tag : tag_78; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1104 = 8'h4f == req_index ? req_tag : tag_79; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1105 = 8'h50 == req_index ? req_tag : tag_80; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1106 = 8'h51 == req_index ? req_tag : tag_81; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1107 = 8'h52 == req_index ? req_tag : tag_82; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1108 = 8'h53 == req_index ? req_tag : tag_83; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1109 = 8'h54 == req_index ? req_tag : tag_84; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1110 = 8'h55 == req_index ? req_tag : tag_85; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1111 = 8'h56 == req_index ? req_tag : tag_86; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1112 = 8'h57 == req_index ? req_tag : tag_87; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1113 = 8'h58 == req_index ? req_tag : tag_88; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1114 = 8'h59 == req_index ? req_tag : tag_89; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1115 = 8'h5a == req_index ? req_tag : tag_90; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1116 = 8'h5b == req_index ? req_tag : tag_91; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1117 = 8'h5c == req_index ? req_tag : tag_92; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1118 = 8'h5d == req_index ? req_tag : tag_93; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1119 = 8'h5e == req_index ? req_tag : tag_94; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1120 = 8'h5f == req_index ? req_tag : tag_95; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1121 = 8'h60 == req_index ? req_tag : tag_96; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1122 = 8'h61 == req_index ? req_tag : tag_97; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1123 = 8'h62 == req_index ? req_tag : tag_98; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1124 = 8'h63 == req_index ? req_tag : tag_99; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1125 = 8'h64 == req_index ? req_tag : tag_100; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1126 = 8'h65 == req_index ? req_tag : tag_101; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1127 = 8'h66 == req_index ? req_tag : tag_102; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1128 = 8'h67 == req_index ? req_tag : tag_103; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1129 = 8'h68 == req_index ? req_tag : tag_104; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1130 = 8'h69 == req_index ? req_tag : tag_105; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1131 = 8'h6a == req_index ? req_tag : tag_106; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1132 = 8'h6b == req_index ? req_tag : tag_107; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1133 = 8'h6c == req_index ? req_tag : tag_108; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1134 = 8'h6d == req_index ? req_tag : tag_109; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1135 = 8'h6e == req_index ? req_tag : tag_110; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1136 = 8'h6f == req_index ? req_tag : tag_111; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1137 = 8'h70 == req_index ? req_tag : tag_112; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1138 = 8'h71 == req_index ? req_tag : tag_113; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1139 = 8'h72 == req_index ? req_tag : tag_114; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1140 = 8'h73 == req_index ? req_tag : tag_115; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1141 = 8'h74 == req_index ? req_tag : tag_116; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1142 = 8'h75 == req_index ? req_tag : tag_117; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1143 = 8'h76 == req_index ? req_tag : tag_118; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1144 = 8'h77 == req_index ? req_tag : tag_119; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1145 = 8'h78 == req_index ? req_tag : tag_120; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1146 = 8'h79 == req_index ? req_tag : tag_121; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1147 = 8'h7a == req_index ? req_tag : tag_122; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1148 = 8'h7b == req_index ? req_tag : tag_123; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1149 = 8'h7c == req_index ? req_tag : tag_124; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1150 = 8'h7d == req_index ? req_tag : tag_125; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1151 = 8'h7e == req_index ? req_tag : tag_126; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1152 = 8'h7f == req_index ? req_tag : tag_127; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1153 = 8'h80 == req_index ? req_tag : tag_128; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1154 = 8'h81 == req_index ? req_tag : tag_129; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1155 = 8'h82 == req_index ? req_tag : tag_130; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1156 = 8'h83 == req_index ? req_tag : tag_131; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1157 = 8'h84 == req_index ? req_tag : tag_132; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1158 = 8'h85 == req_index ? req_tag : tag_133; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1159 = 8'h86 == req_index ? req_tag : tag_134; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1160 = 8'h87 == req_index ? req_tag : tag_135; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1161 = 8'h88 == req_index ? req_tag : tag_136; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1162 = 8'h89 == req_index ? req_tag : tag_137; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1163 = 8'h8a == req_index ? req_tag : tag_138; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1164 = 8'h8b == req_index ? req_tag : tag_139; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1165 = 8'h8c == req_index ? req_tag : tag_140; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1166 = 8'h8d == req_index ? req_tag : tag_141; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1167 = 8'h8e == req_index ? req_tag : tag_142; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1168 = 8'h8f == req_index ? req_tag : tag_143; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1169 = 8'h90 == req_index ? req_tag : tag_144; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1170 = 8'h91 == req_index ? req_tag : tag_145; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1171 = 8'h92 == req_index ? req_tag : tag_146; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1172 = 8'h93 == req_index ? req_tag : tag_147; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1173 = 8'h94 == req_index ? req_tag : tag_148; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1174 = 8'h95 == req_index ? req_tag : tag_149; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1175 = 8'h96 == req_index ? req_tag : tag_150; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1176 = 8'h97 == req_index ? req_tag : tag_151; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1177 = 8'h98 == req_index ? req_tag : tag_152; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1178 = 8'h99 == req_index ? req_tag : tag_153; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1179 = 8'h9a == req_index ? req_tag : tag_154; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1180 = 8'h9b == req_index ? req_tag : tag_155; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1181 = 8'h9c == req_index ? req_tag : tag_156; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1182 = 8'h9d == req_index ? req_tag : tag_157; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1183 = 8'h9e == req_index ? req_tag : tag_158; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1184 = 8'h9f == req_index ? req_tag : tag_159; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1185 = 8'ha0 == req_index ? req_tag : tag_160; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1186 = 8'ha1 == req_index ? req_tag : tag_161; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1187 = 8'ha2 == req_index ? req_tag : tag_162; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1188 = 8'ha3 == req_index ? req_tag : tag_163; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1189 = 8'ha4 == req_index ? req_tag : tag_164; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1190 = 8'ha5 == req_index ? req_tag : tag_165; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1191 = 8'ha6 == req_index ? req_tag : tag_166; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1192 = 8'ha7 == req_index ? req_tag : tag_167; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1193 = 8'ha8 == req_index ? req_tag : tag_168; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1194 = 8'ha9 == req_index ? req_tag : tag_169; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1195 = 8'haa == req_index ? req_tag : tag_170; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1196 = 8'hab == req_index ? req_tag : tag_171; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1197 = 8'hac == req_index ? req_tag : tag_172; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1198 = 8'had == req_index ? req_tag : tag_173; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1199 = 8'hae == req_index ? req_tag : tag_174; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1200 = 8'haf == req_index ? req_tag : tag_175; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1201 = 8'hb0 == req_index ? req_tag : tag_176; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1202 = 8'hb1 == req_index ? req_tag : tag_177; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1203 = 8'hb2 == req_index ? req_tag : tag_178; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1204 = 8'hb3 == req_index ? req_tag : tag_179; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1205 = 8'hb4 == req_index ? req_tag : tag_180; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1206 = 8'hb5 == req_index ? req_tag : tag_181; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1207 = 8'hb6 == req_index ? req_tag : tag_182; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1208 = 8'hb7 == req_index ? req_tag : tag_183; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1209 = 8'hb8 == req_index ? req_tag : tag_184; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1210 = 8'hb9 == req_index ? req_tag : tag_185; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1211 = 8'hba == req_index ? req_tag : tag_186; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1212 = 8'hbb == req_index ? req_tag : tag_187; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1213 = 8'hbc == req_index ? req_tag : tag_188; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1214 = 8'hbd == req_index ? req_tag : tag_189; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1215 = 8'hbe == req_index ? req_tag : tag_190; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1216 = 8'hbf == req_index ? req_tag : tag_191; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1217 = 8'hc0 == req_index ? req_tag : tag_192; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1218 = 8'hc1 == req_index ? req_tag : tag_193; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1219 = 8'hc2 == req_index ? req_tag : tag_194; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1220 = 8'hc3 == req_index ? req_tag : tag_195; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1221 = 8'hc4 == req_index ? req_tag : tag_196; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1222 = 8'hc5 == req_index ? req_tag : tag_197; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1223 = 8'hc6 == req_index ? req_tag : tag_198; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1224 = 8'hc7 == req_index ? req_tag : tag_199; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1225 = 8'hc8 == req_index ? req_tag : tag_200; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1226 = 8'hc9 == req_index ? req_tag : tag_201; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1227 = 8'hca == req_index ? req_tag : tag_202; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1228 = 8'hcb == req_index ? req_tag : tag_203; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1229 = 8'hcc == req_index ? req_tag : tag_204; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1230 = 8'hcd == req_index ? req_tag : tag_205; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1231 = 8'hce == req_index ? req_tag : tag_206; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1232 = 8'hcf == req_index ? req_tag : tag_207; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1233 = 8'hd0 == req_index ? req_tag : tag_208; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1234 = 8'hd1 == req_index ? req_tag : tag_209; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1235 = 8'hd2 == req_index ? req_tag : tag_210; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1236 = 8'hd3 == req_index ? req_tag : tag_211; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1237 = 8'hd4 == req_index ? req_tag : tag_212; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1238 = 8'hd5 == req_index ? req_tag : tag_213; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1239 = 8'hd6 == req_index ? req_tag : tag_214; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1240 = 8'hd7 == req_index ? req_tag : tag_215; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1241 = 8'hd8 == req_index ? req_tag : tag_216; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1242 = 8'hd9 == req_index ? req_tag : tag_217; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1243 = 8'hda == req_index ? req_tag : tag_218; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1244 = 8'hdb == req_index ? req_tag : tag_219; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1245 = 8'hdc == req_index ? req_tag : tag_220; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1246 = 8'hdd == req_index ? req_tag : tag_221; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1247 = 8'hde == req_index ? req_tag : tag_222; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1248 = 8'hdf == req_index ? req_tag : tag_223; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1249 = 8'he0 == req_index ? req_tag : tag_224; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1250 = 8'he1 == req_index ? req_tag : tag_225; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1251 = 8'he2 == req_index ? req_tag : tag_226; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1252 = 8'he3 == req_index ? req_tag : tag_227; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1253 = 8'he4 == req_index ? req_tag : tag_228; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1254 = 8'he5 == req_index ? req_tag : tag_229; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1255 = 8'he6 == req_index ? req_tag : tag_230; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1256 = 8'he7 == req_index ? req_tag : tag_231; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1257 = 8'he8 == req_index ? req_tag : tag_232; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1258 = 8'he9 == req_index ? req_tag : tag_233; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1259 = 8'hea == req_index ? req_tag : tag_234; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1260 = 8'heb == req_index ? req_tag : tag_235; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1261 = 8'hec == req_index ? req_tag : tag_236; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1262 = 8'hed == req_index ? req_tag : tag_237; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1263 = 8'hee == req_index ? req_tag : tag_238; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1264 = 8'hef == req_index ? req_tag : tag_239; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1265 = 8'hf0 == req_index ? req_tag : tag_240; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1266 = 8'hf1 == req_index ? req_tag : tag_241; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1267 = 8'hf2 == req_index ? req_tag : tag_242; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1268 = 8'hf3 == req_index ? req_tag : tag_243; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1269 = 8'hf4 == req_index ? req_tag : tag_244; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1270 = 8'hf5 == req_index ? req_tag : tag_245; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1271 = 8'hf6 == req_index ? req_tag : tag_246; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1272 = 8'hf7 == req_index ? req_tag : tag_247; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1273 = 8'hf8 == req_index ? req_tag : tag_248; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1274 = 8'hf9 == req_index ? req_tag : tag_249; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1275 = 8'hfa == req_index ? req_tag : tag_250; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1276 = 8'hfb == req_index ? req_tag : tag_251; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1277 = 8'hfc == req_index ? req_tag : tag_252; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1278 = 8'hfd == req_index ? req_tag : tag_253; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1279 = 8'hfe == req_index ? req_tag : tag_254; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1280 = 8'hff == req_index ? req_tag : tag_255; // @[Dcache.scala 136:27 Dcache.scala 136:27 Dcache.scala 16:24]
  wire [3:0] _GEN_1281 = 8'h0 == req_index ? req_offset : offset_0; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1282 = 8'h1 == req_index ? req_offset : offset_1; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1283 = 8'h2 == req_index ? req_offset : offset_2; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1284 = 8'h3 == req_index ? req_offset : offset_3; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1285 = 8'h4 == req_index ? req_offset : offset_4; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1286 = 8'h5 == req_index ? req_offset : offset_5; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1287 = 8'h6 == req_index ? req_offset : offset_6; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1288 = 8'h7 == req_index ? req_offset : offset_7; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1289 = 8'h8 == req_index ? req_offset : offset_8; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1290 = 8'h9 == req_index ? req_offset : offset_9; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1291 = 8'ha == req_index ? req_offset : offset_10; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1292 = 8'hb == req_index ? req_offset : offset_11; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1293 = 8'hc == req_index ? req_offset : offset_12; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1294 = 8'hd == req_index ? req_offset : offset_13; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1295 = 8'he == req_index ? req_offset : offset_14; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1296 = 8'hf == req_index ? req_offset : offset_15; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1297 = 8'h10 == req_index ? req_offset : offset_16; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1298 = 8'h11 == req_index ? req_offset : offset_17; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1299 = 8'h12 == req_index ? req_offset : offset_18; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1300 = 8'h13 == req_index ? req_offset : offset_19; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1301 = 8'h14 == req_index ? req_offset : offset_20; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1302 = 8'h15 == req_index ? req_offset : offset_21; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1303 = 8'h16 == req_index ? req_offset : offset_22; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1304 = 8'h17 == req_index ? req_offset : offset_23; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1305 = 8'h18 == req_index ? req_offset : offset_24; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1306 = 8'h19 == req_index ? req_offset : offset_25; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1307 = 8'h1a == req_index ? req_offset : offset_26; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1308 = 8'h1b == req_index ? req_offset : offset_27; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1309 = 8'h1c == req_index ? req_offset : offset_28; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1310 = 8'h1d == req_index ? req_offset : offset_29; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1311 = 8'h1e == req_index ? req_offset : offset_30; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1312 = 8'h1f == req_index ? req_offset : offset_31; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1313 = 8'h20 == req_index ? req_offset : offset_32; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1314 = 8'h21 == req_index ? req_offset : offset_33; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1315 = 8'h22 == req_index ? req_offset : offset_34; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1316 = 8'h23 == req_index ? req_offset : offset_35; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1317 = 8'h24 == req_index ? req_offset : offset_36; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1318 = 8'h25 == req_index ? req_offset : offset_37; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1319 = 8'h26 == req_index ? req_offset : offset_38; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1320 = 8'h27 == req_index ? req_offset : offset_39; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1321 = 8'h28 == req_index ? req_offset : offset_40; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1322 = 8'h29 == req_index ? req_offset : offset_41; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1323 = 8'h2a == req_index ? req_offset : offset_42; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1324 = 8'h2b == req_index ? req_offset : offset_43; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1325 = 8'h2c == req_index ? req_offset : offset_44; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1326 = 8'h2d == req_index ? req_offset : offset_45; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1327 = 8'h2e == req_index ? req_offset : offset_46; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1328 = 8'h2f == req_index ? req_offset : offset_47; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1329 = 8'h30 == req_index ? req_offset : offset_48; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1330 = 8'h31 == req_index ? req_offset : offset_49; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1331 = 8'h32 == req_index ? req_offset : offset_50; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1332 = 8'h33 == req_index ? req_offset : offset_51; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1333 = 8'h34 == req_index ? req_offset : offset_52; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1334 = 8'h35 == req_index ? req_offset : offset_53; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1335 = 8'h36 == req_index ? req_offset : offset_54; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1336 = 8'h37 == req_index ? req_offset : offset_55; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1337 = 8'h38 == req_index ? req_offset : offset_56; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1338 = 8'h39 == req_index ? req_offset : offset_57; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1339 = 8'h3a == req_index ? req_offset : offset_58; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1340 = 8'h3b == req_index ? req_offset : offset_59; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1341 = 8'h3c == req_index ? req_offset : offset_60; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1342 = 8'h3d == req_index ? req_offset : offset_61; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1343 = 8'h3e == req_index ? req_offset : offset_62; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1344 = 8'h3f == req_index ? req_offset : offset_63; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1345 = 8'h40 == req_index ? req_offset : offset_64; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1346 = 8'h41 == req_index ? req_offset : offset_65; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1347 = 8'h42 == req_index ? req_offset : offset_66; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1348 = 8'h43 == req_index ? req_offset : offset_67; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1349 = 8'h44 == req_index ? req_offset : offset_68; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1350 = 8'h45 == req_index ? req_offset : offset_69; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1351 = 8'h46 == req_index ? req_offset : offset_70; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1352 = 8'h47 == req_index ? req_offset : offset_71; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1353 = 8'h48 == req_index ? req_offset : offset_72; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1354 = 8'h49 == req_index ? req_offset : offset_73; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1355 = 8'h4a == req_index ? req_offset : offset_74; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1356 = 8'h4b == req_index ? req_offset : offset_75; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1357 = 8'h4c == req_index ? req_offset : offset_76; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1358 = 8'h4d == req_index ? req_offset : offset_77; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1359 = 8'h4e == req_index ? req_offset : offset_78; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1360 = 8'h4f == req_index ? req_offset : offset_79; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1361 = 8'h50 == req_index ? req_offset : offset_80; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1362 = 8'h51 == req_index ? req_offset : offset_81; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1363 = 8'h52 == req_index ? req_offset : offset_82; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1364 = 8'h53 == req_index ? req_offset : offset_83; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1365 = 8'h54 == req_index ? req_offset : offset_84; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1366 = 8'h55 == req_index ? req_offset : offset_85; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1367 = 8'h56 == req_index ? req_offset : offset_86; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1368 = 8'h57 == req_index ? req_offset : offset_87; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1369 = 8'h58 == req_index ? req_offset : offset_88; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1370 = 8'h59 == req_index ? req_offset : offset_89; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1371 = 8'h5a == req_index ? req_offset : offset_90; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1372 = 8'h5b == req_index ? req_offset : offset_91; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1373 = 8'h5c == req_index ? req_offset : offset_92; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1374 = 8'h5d == req_index ? req_offset : offset_93; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1375 = 8'h5e == req_index ? req_offset : offset_94; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1376 = 8'h5f == req_index ? req_offset : offset_95; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1377 = 8'h60 == req_index ? req_offset : offset_96; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1378 = 8'h61 == req_index ? req_offset : offset_97; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1379 = 8'h62 == req_index ? req_offset : offset_98; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1380 = 8'h63 == req_index ? req_offset : offset_99; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1381 = 8'h64 == req_index ? req_offset : offset_100; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1382 = 8'h65 == req_index ? req_offset : offset_101; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1383 = 8'h66 == req_index ? req_offset : offset_102; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1384 = 8'h67 == req_index ? req_offset : offset_103; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1385 = 8'h68 == req_index ? req_offset : offset_104; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1386 = 8'h69 == req_index ? req_offset : offset_105; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1387 = 8'h6a == req_index ? req_offset : offset_106; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1388 = 8'h6b == req_index ? req_offset : offset_107; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1389 = 8'h6c == req_index ? req_offset : offset_108; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1390 = 8'h6d == req_index ? req_offset : offset_109; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1391 = 8'h6e == req_index ? req_offset : offset_110; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1392 = 8'h6f == req_index ? req_offset : offset_111; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1393 = 8'h70 == req_index ? req_offset : offset_112; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1394 = 8'h71 == req_index ? req_offset : offset_113; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1395 = 8'h72 == req_index ? req_offset : offset_114; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1396 = 8'h73 == req_index ? req_offset : offset_115; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1397 = 8'h74 == req_index ? req_offset : offset_116; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1398 = 8'h75 == req_index ? req_offset : offset_117; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1399 = 8'h76 == req_index ? req_offset : offset_118; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1400 = 8'h77 == req_index ? req_offset : offset_119; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1401 = 8'h78 == req_index ? req_offset : offset_120; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1402 = 8'h79 == req_index ? req_offset : offset_121; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1403 = 8'h7a == req_index ? req_offset : offset_122; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1404 = 8'h7b == req_index ? req_offset : offset_123; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1405 = 8'h7c == req_index ? req_offset : offset_124; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1406 = 8'h7d == req_index ? req_offset : offset_125; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1407 = 8'h7e == req_index ? req_offset : offset_126; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1408 = 8'h7f == req_index ? req_offset : offset_127; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1409 = 8'h80 == req_index ? req_offset : offset_128; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1410 = 8'h81 == req_index ? req_offset : offset_129; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1411 = 8'h82 == req_index ? req_offset : offset_130; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1412 = 8'h83 == req_index ? req_offset : offset_131; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1413 = 8'h84 == req_index ? req_offset : offset_132; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1414 = 8'h85 == req_index ? req_offset : offset_133; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1415 = 8'h86 == req_index ? req_offset : offset_134; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1416 = 8'h87 == req_index ? req_offset : offset_135; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1417 = 8'h88 == req_index ? req_offset : offset_136; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1418 = 8'h89 == req_index ? req_offset : offset_137; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1419 = 8'h8a == req_index ? req_offset : offset_138; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1420 = 8'h8b == req_index ? req_offset : offset_139; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1421 = 8'h8c == req_index ? req_offset : offset_140; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1422 = 8'h8d == req_index ? req_offset : offset_141; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1423 = 8'h8e == req_index ? req_offset : offset_142; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1424 = 8'h8f == req_index ? req_offset : offset_143; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1425 = 8'h90 == req_index ? req_offset : offset_144; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1426 = 8'h91 == req_index ? req_offset : offset_145; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1427 = 8'h92 == req_index ? req_offset : offset_146; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1428 = 8'h93 == req_index ? req_offset : offset_147; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1429 = 8'h94 == req_index ? req_offset : offset_148; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1430 = 8'h95 == req_index ? req_offset : offset_149; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1431 = 8'h96 == req_index ? req_offset : offset_150; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1432 = 8'h97 == req_index ? req_offset : offset_151; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1433 = 8'h98 == req_index ? req_offset : offset_152; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1434 = 8'h99 == req_index ? req_offset : offset_153; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1435 = 8'h9a == req_index ? req_offset : offset_154; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1436 = 8'h9b == req_index ? req_offset : offset_155; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1437 = 8'h9c == req_index ? req_offset : offset_156; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1438 = 8'h9d == req_index ? req_offset : offset_157; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1439 = 8'h9e == req_index ? req_offset : offset_158; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1440 = 8'h9f == req_index ? req_offset : offset_159; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1441 = 8'ha0 == req_index ? req_offset : offset_160; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1442 = 8'ha1 == req_index ? req_offset : offset_161; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1443 = 8'ha2 == req_index ? req_offset : offset_162; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1444 = 8'ha3 == req_index ? req_offset : offset_163; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1445 = 8'ha4 == req_index ? req_offset : offset_164; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1446 = 8'ha5 == req_index ? req_offset : offset_165; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1447 = 8'ha6 == req_index ? req_offset : offset_166; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1448 = 8'ha7 == req_index ? req_offset : offset_167; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1449 = 8'ha8 == req_index ? req_offset : offset_168; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1450 = 8'ha9 == req_index ? req_offset : offset_169; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1451 = 8'haa == req_index ? req_offset : offset_170; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1452 = 8'hab == req_index ? req_offset : offset_171; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1453 = 8'hac == req_index ? req_offset : offset_172; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1454 = 8'had == req_index ? req_offset : offset_173; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1455 = 8'hae == req_index ? req_offset : offset_174; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1456 = 8'haf == req_index ? req_offset : offset_175; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1457 = 8'hb0 == req_index ? req_offset : offset_176; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1458 = 8'hb1 == req_index ? req_offset : offset_177; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1459 = 8'hb2 == req_index ? req_offset : offset_178; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1460 = 8'hb3 == req_index ? req_offset : offset_179; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1461 = 8'hb4 == req_index ? req_offset : offset_180; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1462 = 8'hb5 == req_index ? req_offset : offset_181; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1463 = 8'hb6 == req_index ? req_offset : offset_182; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1464 = 8'hb7 == req_index ? req_offset : offset_183; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1465 = 8'hb8 == req_index ? req_offset : offset_184; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1466 = 8'hb9 == req_index ? req_offset : offset_185; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1467 = 8'hba == req_index ? req_offset : offset_186; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1468 = 8'hbb == req_index ? req_offset : offset_187; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1469 = 8'hbc == req_index ? req_offset : offset_188; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1470 = 8'hbd == req_index ? req_offset : offset_189; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1471 = 8'hbe == req_index ? req_offset : offset_190; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1472 = 8'hbf == req_index ? req_offset : offset_191; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1473 = 8'hc0 == req_index ? req_offset : offset_192; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1474 = 8'hc1 == req_index ? req_offset : offset_193; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1475 = 8'hc2 == req_index ? req_offset : offset_194; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1476 = 8'hc3 == req_index ? req_offset : offset_195; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1477 = 8'hc4 == req_index ? req_offset : offset_196; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1478 = 8'hc5 == req_index ? req_offset : offset_197; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1479 = 8'hc6 == req_index ? req_offset : offset_198; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1480 = 8'hc7 == req_index ? req_offset : offset_199; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1481 = 8'hc8 == req_index ? req_offset : offset_200; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1482 = 8'hc9 == req_index ? req_offset : offset_201; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1483 = 8'hca == req_index ? req_offset : offset_202; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1484 = 8'hcb == req_index ? req_offset : offset_203; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1485 = 8'hcc == req_index ? req_offset : offset_204; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1486 = 8'hcd == req_index ? req_offset : offset_205; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1487 = 8'hce == req_index ? req_offset : offset_206; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1488 = 8'hcf == req_index ? req_offset : offset_207; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1489 = 8'hd0 == req_index ? req_offset : offset_208; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1490 = 8'hd1 == req_index ? req_offset : offset_209; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1491 = 8'hd2 == req_index ? req_offset : offset_210; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1492 = 8'hd3 == req_index ? req_offset : offset_211; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1493 = 8'hd4 == req_index ? req_offset : offset_212; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1494 = 8'hd5 == req_index ? req_offset : offset_213; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1495 = 8'hd6 == req_index ? req_offset : offset_214; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1496 = 8'hd7 == req_index ? req_offset : offset_215; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1497 = 8'hd8 == req_index ? req_offset : offset_216; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1498 = 8'hd9 == req_index ? req_offset : offset_217; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1499 = 8'hda == req_index ? req_offset : offset_218; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1500 = 8'hdb == req_index ? req_offset : offset_219; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1501 = 8'hdc == req_index ? req_offset : offset_220; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1502 = 8'hdd == req_index ? req_offset : offset_221; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1503 = 8'hde == req_index ? req_offset : offset_222; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1504 = 8'hdf == req_index ? req_offset : offset_223; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1505 = 8'he0 == req_index ? req_offset : offset_224; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1506 = 8'he1 == req_index ? req_offset : offset_225; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1507 = 8'he2 == req_index ? req_offset : offset_226; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1508 = 8'he3 == req_index ? req_offset : offset_227; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1509 = 8'he4 == req_index ? req_offset : offset_228; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1510 = 8'he5 == req_index ? req_offset : offset_229; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1511 = 8'he6 == req_index ? req_offset : offset_230; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1512 = 8'he7 == req_index ? req_offset : offset_231; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1513 = 8'he8 == req_index ? req_offset : offset_232; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1514 = 8'he9 == req_index ? req_offset : offset_233; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1515 = 8'hea == req_index ? req_offset : offset_234; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1516 = 8'heb == req_index ? req_offset : offset_235; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1517 = 8'hec == req_index ? req_offset : offset_236; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1518 = 8'hed == req_index ? req_offset : offset_237; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1519 = 8'hee == req_index ? req_offset : offset_238; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1520 = 8'hef == req_index ? req_offset : offset_239; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1521 = 8'hf0 == req_index ? req_offset : offset_240; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1522 = 8'hf1 == req_index ? req_offset : offset_241; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1523 = 8'hf2 == req_index ? req_offset : offset_242; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1524 = 8'hf3 == req_index ? req_offset : offset_243; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1525 = 8'hf4 == req_index ? req_offset : offset_244; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1526 = 8'hf5 == req_index ? req_offset : offset_245; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1527 = 8'hf6 == req_index ? req_offset : offset_246; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1528 = 8'hf7 == req_index ? req_offset : offset_247; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1529 = 8'hf8 == req_index ? req_offset : offset_248; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1530 = 8'hf9 == req_index ? req_offset : offset_249; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1531 = 8'hfa == req_index ? req_offset : offset_250; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1532 = 8'hfb == req_index ? req_offset : offset_251; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1533 = 8'hfc == req_index ? req_offset : offset_252; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1534 = 8'hfd == req_index ? req_offset : offset_253; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1535 = 8'hfe == req_index ? req_offset : offset_254; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1536 = 8'hff == req_index ? req_offset : offset_255; // @[Dcache.scala 137:27 Dcache.scala 137:27 Dcache.scala 19:24]
  wire [127:0] _cache_wdata_T_1 = {valid_wdata,64'h0}; // @[Cat.scala 30:58]
  wire [127:0] _cache_wdata_T_2 = {64'h0,valid_wdata}; // @[Cat.scala 30:58]
  wire [127:0] _cache_wdata_T_3 = req_offset[3] ? _cache_wdata_T_1 : _cache_wdata_T_2; // @[Dcache.scala 140:33]
  wire [127:0] _cache_strb_T_1 = {valid_strb,64'h0}; // @[Cat.scala 30:58]
  wire [127:0] _cache_strb_T_2 = {64'h0,valid_strb}; // @[Cat.scala 30:58]
  wire [127:0] _cache_strb_T_3 = req_offset[3] ? _cache_strb_T_1 : _cache_strb_T_2; // @[Dcache.scala 141:33]
  wire  _GEN_1537 = 8'h0 == req_index ? io_dmem_data_req : dirty_0; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1538 = 8'h1 == req_index ? io_dmem_data_req : dirty_1; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1539 = 8'h2 == req_index ? io_dmem_data_req : dirty_2; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1540 = 8'h3 == req_index ? io_dmem_data_req : dirty_3; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1541 = 8'h4 == req_index ? io_dmem_data_req : dirty_4; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1542 = 8'h5 == req_index ? io_dmem_data_req : dirty_5; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1543 = 8'h6 == req_index ? io_dmem_data_req : dirty_6; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1544 = 8'h7 == req_index ? io_dmem_data_req : dirty_7; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1545 = 8'h8 == req_index ? io_dmem_data_req : dirty_8; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1546 = 8'h9 == req_index ? io_dmem_data_req : dirty_9; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1547 = 8'ha == req_index ? io_dmem_data_req : dirty_10; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1548 = 8'hb == req_index ? io_dmem_data_req : dirty_11; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1549 = 8'hc == req_index ? io_dmem_data_req : dirty_12; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1550 = 8'hd == req_index ? io_dmem_data_req : dirty_13; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1551 = 8'he == req_index ? io_dmem_data_req : dirty_14; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1552 = 8'hf == req_index ? io_dmem_data_req : dirty_15; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1553 = 8'h10 == req_index ? io_dmem_data_req : dirty_16; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1554 = 8'h11 == req_index ? io_dmem_data_req : dirty_17; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1555 = 8'h12 == req_index ? io_dmem_data_req : dirty_18; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1556 = 8'h13 == req_index ? io_dmem_data_req : dirty_19; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1557 = 8'h14 == req_index ? io_dmem_data_req : dirty_20; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1558 = 8'h15 == req_index ? io_dmem_data_req : dirty_21; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1559 = 8'h16 == req_index ? io_dmem_data_req : dirty_22; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1560 = 8'h17 == req_index ? io_dmem_data_req : dirty_23; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1561 = 8'h18 == req_index ? io_dmem_data_req : dirty_24; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1562 = 8'h19 == req_index ? io_dmem_data_req : dirty_25; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1563 = 8'h1a == req_index ? io_dmem_data_req : dirty_26; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1564 = 8'h1b == req_index ? io_dmem_data_req : dirty_27; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1565 = 8'h1c == req_index ? io_dmem_data_req : dirty_28; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1566 = 8'h1d == req_index ? io_dmem_data_req : dirty_29; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1567 = 8'h1e == req_index ? io_dmem_data_req : dirty_30; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1568 = 8'h1f == req_index ? io_dmem_data_req : dirty_31; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1569 = 8'h20 == req_index ? io_dmem_data_req : dirty_32; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1570 = 8'h21 == req_index ? io_dmem_data_req : dirty_33; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1571 = 8'h22 == req_index ? io_dmem_data_req : dirty_34; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1572 = 8'h23 == req_index ? io_dmem_data_req : dirty_35; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1573 = 8'h24 == req_index ? io_dmem_data_req : dirty_36; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1574 = 8'h25 == req_index ? io_dmem_data_req : dirty_37; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1575 = 8'h26 == req_index ? io_dmem_data_req : dirty_38; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1576 = 8'h27 == req_index ? io_dmem_data_req : dirty_39; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1577 = 8'h28 == req_index ? io_dmem_data_req : dirty_40; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1578 = 8'h29 == req_index ? io_dmem_data_req : dirty_41; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1579 = 8'h2a == req_index ? io_dmem_data_req : dirty_42; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1580 = 8'h2b == req_index ? io_dmem_data_req : dirty_43; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1581 = 8'h2c == req_index ? io_dmem_data_req : dirty_44; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1582 = 8'h2d == req_index ? io_dmem_data_req : dirty_45; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1583 = 8'h2e == req_index ? io_dmem_data_req : dirty_46; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1584 = 8'h2f == req_index ? io_dmem_data_req : dirty_47; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1585 = 8'h30 == req_index ? io_dmem_data_req : dirty_48; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1586 = 8'h31 == req_index ? io_dmem_data_req : dirty_49; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1587 = 8'h32 == req_index ? io_dmem_data_req : dirty_50; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1588 = 8'h33 == req_index ? io_dmem_data_req : dirty_51; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1589 = 8'h34 == req_index ? io_dmem_data_req : dirty_52; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1590 = 8'h35 == req_index ? io_dmem_data_req : dirty_53; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1591 = 8'h36 == req_index ? io_dmem_data_req : dirty_54; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1592 = 8'h37 == req_index ? io_dmem_data_req : dirty_55; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1593 = 8'h38 == req_index ? io_dmem_data_req : dirty_56; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1594 = 8'h39 == req_index ? io_dmem_data_req : dirty_57; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1595 = 8'h3a == req_index ? io_dmem_data_req : dirty_58; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1596 = 8'h3b == req_index ? io_dmem_data_req : dirty_59; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1597 = 8'h3c == req_index ? io_dmem_data_req : dirty_60; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1598 = 8'h3d == req_index ? io_dmem_data_req : dirty_61; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1599 = 8'h3e == req_index ? io_dmem_data_req : dirty_62; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1600 = 8'h3f == req_index ? io_dmem_data_req : dirty_63; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1601 = 8'h40 == req_index ? io_dmem_data_req : dirty_64; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1602 = 8'h41 == req_index ? io_dmem_data_req : dirty_65; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1603 = 8'h42 == req_index ? io_dmem_data_req : dirty_66; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1604 = 8'h43 == req_index ? io_dmem_data_req : dirty_67; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1605 = 8'h44 == req_index ? io_dmem_data_req : dirty_68; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1606 = 8'h45 == req_index ? io_dmem_data_req : dirty_69; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1607 = 8'h46 == req_index ? io_dmem_data_req : dirty_70; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1608 = 8'h47 == req_index ? io_dmem_data_req : dirty_71; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1609 = 8'h48 == req_index ? io_dmem_data_req : dirty_72; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1610 = 8'h49 == req_index ? io_dmem_data_req : dirty_73; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1611 = 8'h4a == req_index ? io_dmem_data_req : dirty_74; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1612 = 8'h4b == req_index ? io_dmem_data_req : dirty_75; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1613 = 8'h4c == req_index ? io_dmem_data_req : dirty_76; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1614 = 8'h4d == req_index ? io_dmem_data_req : dirty_77; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1615 = 8'h4e == req_index ? io_dmem_data_req : dirty_78; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1616 = 8'h4f == req_index ? io_dmem_data_req : dirty_79; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1617 = 8'h50 == req_index ? io_dmem_data_req : dirty_80; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1618 = 8'h51 == req_index ? io_dmem_data_req : dirty_81; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1619 = 8'h52 == req_index ? io_dmem_data_req : dirty_82; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1620 = 8'h53 == req_index ? io_dmem_data_req : dirty_83; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1621 = 8'h54 == req_index ? io_dmem_data_req : dirty_84; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1622 = 8'h55 == req_index ? io_dmem_data_req : dirty_85; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1623 = 8'h56 == req_index ? io_dmem_data_req : dirty_86; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1624 = 8'h57 == req_index ? io_dmem_data_req : dirty_87; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1625 = 8'h58 == req_index ? io_dmem_data_req : dirty_88; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1626 = 8'h59 == req_index ? io_dmem_data_req : dirty_89; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1627 = 8'h5a == req_index ? io_dmem_data_req : dirty_90; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1628 = 8'h5b == req_index ? io_dmem_data_req : dirty_91; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1629 = 8'h5c == req_index ? io_dmem_data_req : dirty_92; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1630 = 8'h5d == req_index ? io_dmem_data_req : dirty_93; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1631 = 8'h5e == req_index ? io_dmem_data_req : dirty_94; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1632 = 8'h5f == req_index ? io_dmem_data_req : dirty_95; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1633 = 8'h60 == req_index ? io_dmem_data_req : dirty_96; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1634 = 8'h61 == req_index ? io_dmem_data_req : dirty_97; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1635 = 8'h62 == req_index ? io_dmem_data_req : dirty_98; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1636 = 8'h63 == req_index ? io_dmem_data_req : dirty_99; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1637 = 8'h64 == req_index ? io_dmem_data_req : dirty_100; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1638 = 8'h65 == req_index ? io_dmem_data_req : dirty_101; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1639 = 8'h66 == req_index ? io_dmem_data_req : dirty_102; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1640 = 8'h67 == req_index ? io_dmem_data_req : dirty_103; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1641 = 8'h68 == req_index ? io_dmem_data_req : dirty_104; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1642 = 8'h69 == req_index ? io_dmem_data_req : dirty_105; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1643 = 8'h6a == req_index ? io_dmem_data_req : dirty_106; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1644 = 8'h6b == req_index ? io_dmem_data_req : dirty_107; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1645 = 8'h6c == req_index ? io_dmem_data_req : dirty_108; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1646 = 8'h6d == req_index ? io_dmem_data_req : dirty_109; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1647 = 8'h6e == req_index ? io_dmem_data_req : dirty_110; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1648 = 8'h6f == req_index ? io_dmem_data_req : dirty_111; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1649 = 8'h70 == req_index ? io_dmem_data_req : dirty_112; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1650 = 8'h71 == req_index ? io_dmem_data_req : dirty_113; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1651 = 8'h72 == req_index ? io_dmem_data_req : dirty_114; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1652 = 8'h73 == req_index ? io_dmem_data_req : dirty_115; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1653 = 8'h74 == req_index ? io_dmem_data_req : dirty_116; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1654 = 8'h75 == req_index ? io_dmem_data_req : dirty_117; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1655 = 8'h76 == req_index ? io_dmem_data_req : dirty_118; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1656 = 8'h77 == req_index ? io_dmem_data_req : dirty_119; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1657 = 8'h78 == req_index ? io_dmem_data_req : dirty_120; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1658 = 8'h79 == req_index ? io_dmem_data_req : dirty_121; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1659 = 8'h7a == req_index ? io_dmem_data_req : dirty_122; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1660 = 8'h7b == req_index ? io_dmem_data_req : dirty_123; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1661 = 8'h7c == req_index ? io_dmem_data_req : dirty_124; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1662 = 8'h7d == req_index ? io_dmem_data_req : dirty_125; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1663 = 8'h7e == req_index ? io_dmem_data_req : dirty_126; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1664 = 8'h7f == req_index ? io_dmem_data_req : dirty_127; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1665 = 8'h80 == req_index ? io_dmem_data_req : dirty_128; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1666 = 8'h81 == req_index ? io_dmem_data_req : dirty_129; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1667 = 8'h82 == req_index ? io_dmem_data_req : dirty_130; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1668 = 8'h83 == req_index ? io_dmem_data_req : dirty_131; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1669 = 8'h84 == req_index ? io_dmem_data_req : dirty_132; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1670 = 8'h85 == req_index ? io_dmem_data_req : dirty_133; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1671 = 8'h86 == req_index ? io_dmem_data_req : dirty_134; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1672 = 8'h87 == req_index ? io_dmem_data_req : dirty_135; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1673 = 8'h88 == req_index ? io_dmem_data_req : dirty_136; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1674 = 8'h89 == req_index ? io_dmem_data_req : dirty_137; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1675 = 8'h8a == req_index ? io_dmem_data_req : dirty_138; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1676 = 8'h8b == req_index ? io_dmem_data_req : dirty_139; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1677 = 8'h8c == req_index ? io_dmem_data_req : dirty_140; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1678 = 8'h8d == req_index ? io_dmem_data_req : dirty_141; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1679 = 8'h8e == req_index ? io_dmem_data_req : dirty_142; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1680 = 8'h8f == req_index ? io_dmem_data_req : dirty_143; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1681 = 8'h90 == req_index ? io_dmem_data_req : dirty_144; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1682 = 8'h91 == req_index ? io_dmem_data_req : dirty_145; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1683 = 8'h92 == req_index ? io_dmem_data_req : dirty_146; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1684 = 8'h93 == req_index ? io_dmem_data_req : dirty_147; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1685 = 8'h94 == req_index ? io_dmem_data_req : dirty_148; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1686 = 8'h95 == req_index ? io_dmem_data_req : dirty_149; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1687 = 8'h96 == req_index ? io_dmem_data_req : dirty_150; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1688 = 8'h97 == req_index ? io_dmem_data_req : dirty_151; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1689 = 8'h98 == req_index ? io_dmem_data_req : dirty_152; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1690 = 8'h99 == req_index ? io_dmem_data_req : dirty_153; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1691 = 8'h9a == req_index ? io_dmem_data_req : dirty_154; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1692 = 8'h9b == req_index ? io_dmem_data_req : dirty_155; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1693 = 8'h9c == req_index ? io_dmem_data_req : dirty_156; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1694 = 8'h9d == req_index ? io_dmem_data_req : dirty_157; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1695 = 8'h9e == req_index ? io_dmem_data_req : dirty_158; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1696 = 8'h9f == req_index ? io_dmem_data_req : dirty_159; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1697 = 8'ha0 == req_index ? io_dmem_data_req : dirty_160; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1698 = 8'ha1 == req_index ? io_dmem_data_req : dirty_161; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1699 = 8'ha2 == req_index ? io_dmem_data_req : dirty_162; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1700 = 8'ha3 == req_index ? io_dmem_data_req : dirty_163; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1701 = 8'ha4 == req_index ? io_dmem_data_req : dirty_164; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1702 = 8'ha5 == req_index ? io_dmem_data_req : dirty_165; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1703 = 8'ha6 == req_index ? io_dmem_data_req : dirty_166; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1704 = 8'ha7 == req_index ? io_dmem_data_req : dirty_167; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1705 = 8'ha8 == req_index ? io_dmem_data_req : dirty_168; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1706 = 8'ha9 == req_index ? io_dmem_data_req : dirty_169; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1707 = 8'haa == req_index ? io_dmem_data_req : dirty_170; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1708 = 8'hab == req_index ? io_dmem_data_req : dirty_171; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1709 = 8'hac == req_index ? io_dmem_data_req : dirty_172; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1710 = 8'had == req_index ? io_dmem_data_req : dirty_173; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1711 = 8'hae == req_index ? io_dmem_data_req : dirty_174; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1712 = 8'haf == req_index ? io_dmem_data_req : dirty_175; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1713 = 8'hb0 == req_index ? io_dmem_data_req : dirty_176; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1714 = 8'hb1 == req_index ? io_dmem_data_req : dirty_177; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1715 = 8'hb2 == req_index ? io_dmem_data_req : dirty_178; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1716 = 8'hb3 == req_index ? io_dmem_data_req : dirty_179; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1717 = 8'hb4 == req_index ? io_dmem_data_req : dirty_180; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1718 = 8'hb5 == req_index ? io_dmem_data_req : dirty_181; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1719 = 8'hb6 == req_index ? io_dmem_data_req : dirty_182; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1720 = 8'hb7 == req_index ? io_dmem_data_req : dirty_183; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1721 = 8'hb8 == req_index ? io_dmem_data_req : dirty_184; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1722 = 8'hb9 == req_index ? io_dmem_data_req : dirty_185; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1723 = 8'hba == req_index ? io_dmem_data_req : dirty_186; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1724 = 8'hbb == req_index ? io_dmem_data_req : dirty_187; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1725 = 8'hbc == req_index ? io_dmem_data_req : dirty_188; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1726 = 8'hbd == req_index ? io_dmem_data_req : dirty_189; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1727 = 8'hbe == req_index ? io_dmem_data_req : dirty_190; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1728 = 8'hbf == req_index ? io_dmem_data_req : dirty_191; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1729 = 8'hc0 == req_index ? io_dmem_data_req : dirty_192; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1730 = 8'hc1 == req_index ? io_dmem_data_req : dirty_193; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1731 = 8'hc2 == req_index ? io_dmem_data_req : dirty_194; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1732 = 8'hc3 == req_index ? io_dmem_data_req : dirty_195; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1733 = 8'hc4 == req_index ? io_dmem_data_req : dirty_196; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1734 = 8'hc5 == req_index ? io_dmem_data_req : dirty_197; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1735 = 8'hc6 == req_index ? io_dmem_data_req : dirty_198; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1736 = 8'hc7 == req_index ? io_dmem_data_req : dirty_199; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1737 = 8'hc8 == req_index ? io_dmem_data_req : dirty_200; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1738 = 8'hc9 == req_index ? io_dmem_data_req : dirty_201; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1739 = 8'hca == req_index ? io_dmem_data_req : dirty_202; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1740 = 8'hcb == req_index ? io_dmem_data_req : dirty_203; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1741 = 8'hcc == req_index ? io_dmem_data_req : dirty_204; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1742 = 8'hcd == req_index ? io_dmem_data_req : dirty_205; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1743 = 8'hce == req_index ? io_dmem_data_req : dirty_206; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1744 = 8'hcf == req_index ? io_dmem_data_req : dirty_207; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1745 = 8'hd0 == req_index ? io_dmem_data_req : dirty_208; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1746 = 8'hd1 == req_index ? io_dmem_data_req : dirty_209; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1747 = 8'hd2 == req_index ? io_dmem_data_req : dirty_210; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1748 = 8'hd3 == req_index ? io_dmem_data_req : dirty_211; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1749 = 8'hd4 == req_index ? io_dmem_data_req : dirty_212; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1750 = 8'hd5 == req_index ? io_dmem_data_req : dirty_213; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1751 = 8'hd6 == req_index ? io_dmem_data_req : dirty_214; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1752 = 8'hd7 == req_index ? io_dmem_data_req : dirty_215; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1753 = 8'hd8 == req_index ? io_dmem_data_req : dirty_216; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1754 = 8'hd9 == req_index ? io_dmem_data_req : dirty_217; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1755 = 8'hda == req_index ? io_dmem_data_req : dirty_218; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1756 = 8'hdb == req_index ? io_dmem_data_req : dirty_219; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1757 = 8'hdc == req_index ? io_dmem_data_req : dirty_220; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1758 = 8'hdd == req_index ? io_dmem_data_req : dirty_221; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1759 = 8'hde == req_index ? io_dmem_data_req : dirty_222; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1760 = 8'hdf == req_index ? io_dmem_data_req : dirty_223; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1761 = 8'he0 == req_index ? io_dmem_data_req : dirty_224; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1762 = 8'he1 == req_index ? io_dmem_data_req : dirty_225; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1763 = 8'he2 == req_index ? io_dmem_data_req : dirty_226; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1764 = 8'he3 == req_index ? io_dmem_data_req : dirty_227; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1765 = 8'he4 == req_index ? io_dmem_data_req : dirty_228; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1766 = 8'he5 == req_index ? io_dmem_data_req : dirty_229; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1767 = 8'he6 == req_index ? io_dmem_data_req : dirty_230; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1768 = 8'he7 == req_index ? io_dmem_data_req : dirty_231; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1769 = 8'he8 == req_index ? io_dmem_data_req : dirty_232; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1770 = 8'he9 == req_index ? io_dmem_data_req : dirty_233; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1771 = 8'hea == req_index ? io_dmem_data_req : dirty_234; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1772 = 8'heb == req_index ? io_dmem_data_req : dirty_235; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1773 = 8'hec == req_index ? io_dmem_data_req : dirty_236; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1774 = 8'hed == req_index ? io_dmem_data_req : dirty_237; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1775 = 8'hee == req_index ? io_dmem_data_req : dirty_238; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1776 = 8'hef == req_index ? io_dmem_data_req : dirty_239; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1777 = 8'hf0 == req_index ? io_dmem_data_req : dirty_240; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1778 = 8'hf1 == req_index ? io_dmem_data_req : dirty_241; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1779 = 8'hf2 == req_index ? io_dmem_data_req : dirty_242; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1780 = 8'hf3 == req_index ? io_dmem_data_req : dirty_243; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1781 = 8'hf4 == req_index ? io_dmem_data_req : dirty_244; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1782 = 8'hf5 == req_index ? io_dmem_data_req : dirty_245; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1783 = 8'hf6 == req_index ? io_dmem_data_req : dirty_246; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1784 = 8'hf7 == req_index ? io_dmem_data_req : dirty_247; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1785 = 8'hf8 == req_index ? io_dmem_data_req : dirty_248; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1786 = 8'hf9 == req_index ? io_dmem_data_req : dirty_249; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1787 = 8'hfa == req_index ? io_dmem_data_req : dirty_250; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1788 = 8'hfb == req_index ? io_dmem_data_req : dirty_251; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1789 = 8'hfc == req_index ? io_dmem_data_req : dirty_252; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1790 = 8'hfd == req_index ? io_dmem_data_req : dirty_253; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1791 = 8'hfe == req_index ? io_dmem_data_req : dirty_254; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1792 = 8'hff == req_index ? io_dmem_data_req : dirty_255; // @[Dcache.scala 143:28 Dcache.scala 143:28 Dcache.scala 18:24]
  wire  _GEN_1793 = ~_GEN_767 ? _GEN_1537 : dirty_0; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1794 = ~_GEN_767 ? _GEN_1538 : dirty_1; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1795 = ~_GEN_767 ? _GEN_1539 : dirty_2; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1796 = ~_GEN_767 ? _GEN_1540 : dirty_3; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1797 = ~_GEN_767 ? _GEN_1541 : dirty_4; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1798 = ~_GEN_767 ? _GEN_1542 : dirty_5; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1799 = ~_GEN_767 ? _GEN_1543 : dirty_6; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1800 = ~_GEN_767 ? _GEN_1544 : dirty_7; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1801 = ~_GEN_767 ? _GEN_1545 : dirty_8; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1802 = ~_GEN_767 ? _GEN_1546 : dirty_9; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1803 = ~_GEN_767 ? _GEN_1547 : dirty_10; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1804 = ~_GEN_767 ? _GEN_1548 : dirty_11; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1805 = ~_GEN_767 ? _GEN_1549 : dirty_12; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1806 = ~_GEN_767 ? _GEN_1550 : dirty_13; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1807 = ~_GEN_767 ? _GEN_1551 : dirty_14; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1808 = ~_GEN_767 ? _GEN_1552 : dirty_15; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1809 = ~_GEN_767 ? _GEN_1553 : dirty_16; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1810 = ~_GEN_767 ? _GEN_1554 : dirty_17; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1811 = ~_GEN_767 ? _GEN_1555 : dirty_18; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1812 = ~_GEN_767 ? _GEN_1556 : dirty_19; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1813 = ~_GEN_767 ? _GEN_1557 : dirty_20; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1814 = ~_GEN_767 ? _GEN_1558 : dirty_21; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1815 = ~_GEN_767 ? _GEN_1559 : dirty_22; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1816 = ~_GEN_767 ? _GEN_1560 : dirty_23; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1817 = ~_GEN_767 ? _GEN_1561 : dirty_24; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1818 = ~_GEN_767 ? _GEN_1562 : dirty_25; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1819 = ~_GEN_767 ? _GEN_1563 : dirty_26; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1820 = ~_GEN_767 ? _GEN_1564 : dirty_27; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1821 = ~_GEN_767 ? _GEN_1565 : dirty_28; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1822 = ~_GEN_767 ? _GEN_1566 : dirty_29; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1823 = ~_GEN_767 ? _GEN_1567 : dirty_30; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1824 = ~_GEN_767 ? _GEN_1568 : dirty_31; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1825 = ~_GEN_767 ? _GEN_1569 : dirty_32; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1826 = ~_GEN_767 ? _GEN_1570 : dirty_33; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1827 = ~_GEN_767 ? _GEN_1571 : dirty_34; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1828 = ~_GEN_767 ? _GEN_1572 : dirty_35; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1829 = ~_GEN_767 ? _GEN_1573 : dirty_36; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1830 = ~_GEN_767 ? _GEN_1574 : dirty_37; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1831 = ~_GEN_767 ? _GEN_1575 : dirty_38; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1832 = ~_GEN_767 ? _GEN_1576 : dirty_39; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1833 = ~_GEN_767 ? _GEN_1577 : dirty_40; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1834 = ~_GEN_767 ? _GEN_1578 : dirty_41; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1835 = ~_GEN_767 ? _GEN_1579 : dirty_42; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1836 = ~_GEN_767 ? _GEN_1580 : dirty_43; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1837 = ~_GEN_767 ? _GEN_1581 : dirty_44; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1838 = ~_GEN_767 ? _GEN_1582 : dirty_45; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1839 = ~_GEN_767 ? _GEN_1583 : dirty_46; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1840 = ~_GEN_767 ? _GEN_1584 : dirty_47; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1841 = ~_GEN_767 ? _GEN_1585 : dirty_48; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1842 = ~_GEN_767 ? _GEN_1586 : dirty_49; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1843 = ~_GEN_767 ? _GEN_1587 : dirty_50; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1844 = ~_GEN_767 ? _GEN_1588 : dirty_51; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1845 = ~_GEN_767 ? _GEN_1589 : dirty_52; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1846 = ~_GEN_767 ? _GEN_1590 : dirty_53; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1847 = ~_GEN_767 ? _GEN_1591 : dirty_54; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1848 = ~_GEN_767 ? _GEN_1592 : dirty_55; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1849 = ~_GEN_767 ? _GEN_1593 : dirty_56; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1850 = ~_GEN_767 ? _GEN_1594 : dirty_57; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1851 = ~_GEN_767 ? _GEN_1595 : dirty_58; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1852 = ~_GEN_767 ? _GEN_1596 : dirty_59; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1853 = ~_GEN_767 ? _GEN_1597 : dirty_60; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1854 = ~_GEN_767 ? _GEN_1598 : dirty_61; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1855 = ~_GEN_767 ? _GEN_1599 : dirty_62; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1856 = ~_GEN_767 ? _GEN_1600 : dirty_63; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1857 = ~_GEN_767 ? _GEN_1601 : dirty_64; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1858 = ~_GEN_767 ? _GEN_1602 : dirty_65; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1859 = ~_GEN_767 ? _GEN_1603 : dirty_66; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1860 = ~_GEN_767 ? _GEN_1604 : dirty_67; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1861 = ~_GEN_767 ? _GEN_1605 : dirty_68; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1862 = ~_GEN_767 ? _GEN_1606 : dirty_69; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1863 = ~_GEN_767 ? _GEN_1607 : dirty_70; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1864 = ~_GEN_767 ? _GEN_1608 : dirty_71; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1865 = ~_GEN_767 ? _GEN_1609 : dirty_72; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1866 = ~_GEN_767 ? _GEN_1610 : dirty_73; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1867 = ~_GEN_767 ? _GEN_1611 : dirty_74; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1868 = ~_GEN_767 ? _GEN_1612 : dirty_75; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1869 = ~_GEN_767 ? _GEN_1613 : dirty_76; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1870 = ~_GEN_767 ? _GEN_1614 : dirty_77; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1871 = ~_GEN_767 ? _GEN_1615 : dirty_78; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1872 = ~_GEN_767 ? _GEN_1616 : dirty_79; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1873 = ~_GEN_767 ? _GEN_1617 : dirty_80; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1874 = ~_GEN_767 ? _GEN_1618 : dirty_81; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1875 = ~_GEN_767 ? _GEN_1619 : dirty_82; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1876 = ~_GEN_767 ? _GEN_1620 : dirty_83; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1877 = ~_GEN_767 ? _GEN_1621 : dirty_84; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1878 = ~_GEN_767 ? _GEN_1622 : dirty_85; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1879 = ~_GEN_767 ? _GEN_1623 : dirty_86; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1880 = ~_GEN_767 ? _GEN_1624 : dirty_87; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1881 = ~_GEN_767 ? _GEN_1625 : dirty_88; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1882 = ~_GEN_767 ? _GEN_1626 : dirty_89; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1883 = ~_GEN_767 ? _GEN_1627 : dirty_90; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1884 = ~_GEN_767 ? _GEN_1628 : dirty_91; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1885 = ~_GEN_767 ? _GEN_1629 : dirty_92; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1886 = ~_GEN_767 ? _GEN_1630 : dirty_93; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1887 = ~_GEN_767 ? _GEN_1631 : dirty_94; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1888 = ~_GEN_767 ? _GEN_1632 : dirty_95; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1889 = ~_GEN_767 ? _GEN_1633 : dirty_96; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1890 = ~_GEN_767 ? _GEN_1634 : dirty_97; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1891 = ~_GEN_767 ? _GEN_1635 : dirty_98; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1892 = ~_GEN_767 ? _GEN_1636 : dirty_99; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1893 = ~_GEN_767 ? _GEN_1637 : dirty_100; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1894 = ~_GEN_767 ? _GEN_1638 : dirty_101; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1895 = ~_GEN_767 ? _GEN_1639 : dirty_102; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1896 = ~_GEN_767 ? _GEN_1640 : dirty_103; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1897 = ~_GEN_767 ? _GEN_1641 : dirty_104; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1898 = ~_GEN_767 ? _GEN_1642 : dirty_105; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1899 = ~_GEN_767 ? _GEN_1643 : dirty_106; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1900 = ~_GEN_767 ? _GEN_1644 : dirty_107; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1901 = ~_GEN_767 ? _GEN_1645 : dirty_108; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1902 = ~_GEN_767 ? _GEN_1646 : dirty_109; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1903 = ~_GEN_767 ? _GEN_1647 : dirty_110; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1904 = ~_GEN_767 ? _GEN_1648 : dirty_111; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1905 = ~_GEN_767 ? _GEN_1649 : dirty_112; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1906 = ~_GEN_767 ? _GEN_1650 : dirty_113; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1907 = ~_GEN_767 ? _GEN_1651 : dirty_114; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1908 = ~_GEN_767 ? _GEN_1652 : dirty_115; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1909 = ~_GEN_767 ? _GEN_1653 : dirty_116; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1910 = ~_GEN_767 ? _GEN_1654 : dirty_117; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1911 = ~_GEN_767 ? _GEN_1655 : dirty_118; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1912 = ~_GEN_767 ? _GEN_1656 : dirty_119; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1913 = ~_GEN_767 ? _GEN_1657 : dirty_120; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1914 = ~_GEN_767 ? _GEN_1658 : dirty_121; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1915 = ~_GEN_767 ? _GEN_1659 : dirty_122; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1916 = ~_GEN_767 ? _GEN_1660 : dirty_123; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1917 = ~_GEN_767 ? _GEN_1661 : dirty_124; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1918 = ~_GEN_767 ? _GEN_1662 : dirty_125; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1919 = ~_GEN_767 ? _GEN_1663 : dirty_126; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1920 = ~_GEN_767 ? _GEN_1664 : dirty_127; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1921 = ~_GEN_767 ? _GEN_1665 : dirty_128; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1922 = ~_GEN_767 ? _GEN_1666 : dirty_129; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1923 = ~_GEN_767 ? _GEN_1667 : dirty_130; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1924 = ~_GEN_767 ? _GEN_1668 : dirty_131; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1925 = ~_GEN_767 ? _GEN_1669 : dirty_132; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1926 = ~_GEN_767 ? _GEN_1670 : dirty_133; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1927 = ~_GEN_767 ? _GEN_1671 : dirty_134; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1928 = ~_GEN_767 ? _GEN_1672 : dirty_135; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1929 = ~_GEN_767 ? _GEN_1673 : dirty_136; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1930 = ~_GEN_767 ? _GEN_1674 : dirty_137; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1931 = ~_GEN_767 ? _GEN_1675 : dirty_138; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1932 = ~_GEN_767 ? _GEN_1676 : dirty_139; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1933 = ~_GEN_767 ? _GEN_1677 : dirty_140; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1934 = ~_GEN_767 ? _GEN_1678 : dirty_141; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1935 = ~_GEN_767 ? _GEN_1679 : dirty_142; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1936 = ~_GEN_767 ? _GEN_1680 : dirty_143; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1937 = ~_GEN_767 ? _GEN_1681 : dirty_144; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1938 = ~_GEN_767 ? _GEN_1682 : dirty_145; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1939 = ~_GEN_767 ? _GEN_1683 : dirty_146; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1940 = ~_GEN_767 ? _GEN_1684 : dirty_147; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1941 = ~_GEN_767 ? _GEN_1685 : dirty_148; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1942 = ~_GEN_767 ? _GEN_1686 : dirty_149; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1943 = ~_GEN_767 ? _GEN_1687 : dirty_150; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1944 = ~_GEN_767 ? _GEN_1688 : dirty_151; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1945 = ~_GEN_767 ? _GEN_1689 : dirty_152; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1946 = ~_GEN_767 ? _GEN_1690 : dirty_153; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1947 = ~_GEN_767 ? _GEN_1691 : dirty_154; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1948 = ~_GEN_767 ? _GEN_1692 : dirty_155; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1949 = ~_GEN_767 ? _GEN_1693 : dirty_156; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1950 = ~_GEN_767 ? _GEN_1694 : dirty_157; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1951 = ~_GEN_767 ? _GEN_1695 : dirty_158; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1952 = ~_GEN_767 ? _GEN_1696 : dirty_159; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1953 = ~_GEN_767 ? _GEN_1697 : dirty_160; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1954 = ~_GEN_767 ? _GEN_1698 : dirty_161; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1955 = ~_GEN_767 ? _GEN_1699 : dirty_162; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1956 = ~_GEN_767 ? _GEN_1700 : dirty_163; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1957 = ~_GEN_767 ? _GEN_1701 : dirty_164; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1958 = ~_GEN_767 ? _GEN_1702 : dirty_165; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1959 = ~_GEN_767 ? _GEN_1703 : dirty_166; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1960 = ~_GEN_767 ? _GEN_1704 : dirty_167; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1961 = ~_GEN_767 ? _GEN_1705 : dirty_168; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1962 = ~_GEN_767 ? _GEN_1706 : dirty_169; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1963 = ~_GEN_767 ? _GEN_1707 : dirty_170; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1964 = ~_GEN_767 ? _GEN_1708 : dirty_171; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1965 = ~_GEN_767 ? _GEN_1709 : dirty_172; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1966 = ~_GEN_767 ? _GEN_1710 : dirty_173; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1967 = ~_GEN_767 ? _GEN_1711 : dirty_174; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1968 = ~_GEN_767 ? _GEN_1712 : dirty_175; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1969 = ~_GEN_767 ? _GEN_1713 : dirty_176; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1970 = ~_GEN_767 ? _GEN_1714 : dirty_177; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1971 = ~_GEN_767 ? _GEN_1715 : dirty_178; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1972 = ~_GEN_767 ? _GEN_1716 : dirty_179; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1973 = ~_GEN_767 ? _GEN_1717 : dirty_180; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1974 = ~_GEN_767 ? _GEN_1718 : dirty_181; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1975 = ~_GEN_767 ? _GEN_1719 : dirty_182; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1976 = ~_GEN_767 ? _GEN_1720 : dirty_183; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1977 = ~_GEN_767 ? _GEN_1721 : dirty_184; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1978 = ~_GEN_767 ? _GEN_1722 : dirty_185; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1979 = ~_GEN_767 ? _GEN_1723 : dirty_186; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1980 = ~_GEN_767 ? _GEN_1724 : dirty_187; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1981 = ~_GEN_767 ? _GEN_1725 : dirty_188; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1982 = ~_GEN_767 ? _GEN_1726 : dirty_189; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1983 = ~_GEN_767 ? _GEN_1727 : dirty_190; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1984 = ~_GEN_767 ? _GEN_1728 : dirty_191; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1985 = ~_GEN_767 ? _GEN_1729 : dirty_192; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1986 = ~_GEN_767 ? _GEN_1730 : dirty_193; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1987 = ~_GEN_767 ? _GEN_1731 : dirty_194; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1988 = ~_GEN_767 ? _GEN_1732 : dirty_195; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1989 = ~_GEN_767 ? _GEN_1733 : dirty_196; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1990 = ~_GEN_767 ? _GEN_1734 : dirty_197; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1991 = ~_GEN_767 ? _GEN_1735 : dirty_198; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1992 = ~_GEN_767 ? _GEN_1736 : dirty_199; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1993 = ~_GEN_767 ? _GEN_1737 : dirty_200; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1994 = ~_GEN_767 ? _GEN_1738 : dirty_201; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1995 = ~_GEN_767 ? _GEN_1739 : dirty_202; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1996 = ~_GEN_767 ? _GEN_1740 : dirty_203; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1997 = ~_GEN_767 ? _GEN_1741 : dirty_204; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1998 = ~_GEN_767 ? _GEN_1742 : dirty_205; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_1999 = ~_GEN_767 ? _GEN_1743 : dirty_206; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2000 = ~_GEN_767 ? _GEN_1744 : dirty_207; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2001 = ~_GEN_767 ? _GEN_1745 : dirty_208; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2002 = ~_GEN_767 ? _GEN_1746 : dirty_209; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2003 = ~_GEN_767 ? _GEN_1747 : dirty_210; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2004 = ~_GEN_767 ? _GEN_1748 : dirty_211; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2005 = ~_GEN_767 ? _GEN_1749 : dirty_212; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2006 = ~_GEN_767 ? _GEN_1750 : dirty_213; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2007 = ~_GEN_767 ? _GEN_1751 : dirty_214; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2008 = ~_GEN_767 ? _GEN_1752 : dirty_215; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2009 = ~_GEN_767 ? _GEN_1753 : dirty_216; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2010 = ~_GEN_767 ? _GEN_1754 : dirty_217; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2011 = ~_GEN_767 ? _GEN_1755 : dirty_218; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2012 = ~_GEN_767 ? _GEN_1756 : dirty_219; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2013 = ~_GEN_767 ? _GEN_1757 : dirty_220; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2014 = ~_GEN_767 ? _GEN_1758 : dirty_221; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2015 = ~_GEN_767 ? _GEN_1759 : dirty_222; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2016 = ~_GEN_767 ? _GEN_1760 : dirty_223; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2017 = ~_GEN_767 ? _GEN_1761 : dirty_224; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2018 = ~_GEN_767 ? _GEN_1762 : dirty_225; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2019 = ~_GEN_767 ? _GEN_1763 : dirty_226; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2020 = ~_GEN_767 ? _GEN_1764 : dirty_227; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2021 = ~_GEN_767 ? _GEN_1765 : dirty_228; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2022 = ~_GEN_767 ? _GEN_1766 : dirty_229; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2023 = ~_GEN_767 ? _GEN_1767 : dirty_230; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2024 = ~_GEN_767 ? _GEN_1768 : dirty_231; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2025 = ~_GEN_767 ? _GEN_1769 : dirty_232; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2026 = ~_GEN_767 ? _GEN_1770 : dirty_233; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2027 = ~_GEN_767 ? _GEN_1771 : dirty_234; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2028 = ~_GEN_767 ? _GEN_1772 : dirty_235; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2029 = ~_GEN_767 ? _GEN_1773 : dirty_236; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2030 = ~_GEN_767 ? _GEN_1774 : dirty_237; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2031 = ~_GEN_767 ? _GEN_1775 : dirty_238; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2032 = ~_GEN_767 ? _GEN_1776 : dirty_239; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2033 = ~_GEN_767 ? _GEN_1777 : dirty_240; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2034 = ~_GEN_767 ? _GEN_1778 : dirty_241; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2035 = ~_GEN_767 ? _GEN_1779 : dirty_242; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2036 = ~_GEN_767 ? _GEN_1780 : dirty_243; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2037 = ~_GEN_767 ? _GEN_1781 : dirty_244; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2038 = ~_GEN_767 ? _GEN_1782 : dirty_245; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2039 = ~_GEN_767 ? _GEN_1783 : dirty_246; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2040 = ~_GEN_767 ? _GEN_1784 : dirty_247; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2041 = ~_GEN_767 ? _GEN_1785 : dirty_248; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2042 = ~_GEN_767 ? _GEN_1786 : dirty_249; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2043 = ~_GEN_767 ? _GEN_1787 : dirty_250; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2044 = ~_GEN_767 ? _GEN_1788 : dirty_251; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2045 = ~_GEN_767 ? _GEN_1789 : dirty_252; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2046 = ~_GEN_767 ? _GEN_1790 : dirty_253; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2047 = ~_GEN_767 ? _GEN_1791 : dirty_254; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire  _GEN_2048 = ~_GEN_767 ? _GEN_1792 : dirty_255; // @[Dcache.scala 142:34 Dcache.scala 18:24]
  wire [2:0] _GEN_2049 = cache_dirty ? 3'h2 : 3'h4; // @[Dcache.scala 147:31 Dcache.scala 148:15 Dcache.scala 151:15]
  wire  _GEN_2050 = cache_hit ? _GEN_769 : valid_0; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2051 = cache_hit ? _GEN_770 : valid_1; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2052 = cache_hit ? _GEN_771 : valid_2; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2053 = cache_hit ? _GEN_772 : valid_3; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2054 = cache_hit ? _GEN_773 : valid_4; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2055 = cache_hit ? _GEN_774 : valid_5; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2056 = cache_hit ? _GEN_775 : valid_6; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2057 = cache_hit ? _GEN_776 : valid_7; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2058 = cache_hit ? _GEN_777 : valid_8; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2059 = cache_hit ? _GEN_778 : valid_9; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2060 = cache_hit ? _GEN_779 : valid_10; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2061 = cache_hit ? _GEN_780 : valid_11; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2062 = cache_hit ? _GEN_781 : valid_12; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2063 = cache_hit ? _GEN_782 : valid_13; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2064 = cache_hit ? _GEN_783 : valid_14; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2065 = cache_hit ? _GEN_784 : valid_15; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2066 = cache_hit ? _GEN_785 : valid_16; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2067 = cache_hit ? _GEN_786 : valid_17; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2068 = cache_hit ? _GEN_787 : valid_18; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2069 = cache_hit ? _GEN_788 : valid_19; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2070 = cache_hit ? _GEN_789 : valid_20; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2071 = cache_hit ? _GEN_790 : valid_21; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2072 = cache_hit ? _GEN_791 : valid_22; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2073 = cache_hit ? _GEN_792 : valid_23; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2074 = cache_hit ? _GEN_793 : valid_24; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2075 = cache_hit ? _GEN_794 : valid_25; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2076 = cache_hit ? _GEN_795 : valid_26; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2077 = cache_hit ? _GEN_796 : valid_27; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2078 = cache_hit ? _GEN_797 : valid_28; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2079 = cache_hit ? _GEN_798 : valid_29; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2080 = cache_hit ? _GEN_799 : valid_30; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2081 = cache_hit ? _GEN_800 : valid_31; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2082 = cache_hit ? _GEN_801 : valid_32; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2083 = cache_hit ? _GEN_802 : valid_33; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2084 = cache_hit ? _GEN_803 : valid_34; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2085 = cache_hit ? _GEN_804 : valid_35; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2086 = cache_hit ? _GEN_805 : valid_36; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2087 = cache_hit ? _GEN_806 : valid_37; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2088 = cache_hit ? _GEN_807 : valid_38; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2089 = cache_hit ? _GEN_808 : valid_39; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2090 = cache_hit ? _GEN_809 : valid_40; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2091 = cache_hit ? _GEN_810 : valid_41; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2092 = cache_hit ? _GEN_811 : valid_42; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2093 = cache_hit ? _GEN_812 : valid_43; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2094 = cache_hit ? _GEN_813 : valid_44; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2095 = cache_hit ? _GEN_814 : valid_45; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2096 = cache_hit ? _GEN_815 : valid_46; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2097 = cache_hit ? _GEN_816 : valid_47; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2098 = cache_hit ? _GEN_817 : valid_48; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2099 = cache_hit ? _GEN_818 : valid_49; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2100 = cache_hit ? _GEN_819 : valid_50; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2101 = cache_hit ? _GEN_820 : valid_51; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2102 = cache_hit ? _GEN_821 : valid_52; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2103 = cache_hit ? _GEN_822 : valid_53; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2104 = cache_hit ? _GEN_823 : valid_54; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2105 = cache_hit ? _GEN_824 : valid_55; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2106 = cache_hit ? _GEN_825 : valid_56; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2107 = cache_hit ? _GEN_826 : valid_57; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2108 = cache_hit ? _GEN_827 : valid_58; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2109 = cache_hit ? _GEN_828 : valid_59; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2110 = cache_hit ? _GEN_829 : valid_60; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2111 = cache_hit ? _GEN_830 : valid_61; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2112 = cache_hit ? _GEN_831 : valid_62; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2113 = cache_hit ? _GEN_832 : valid_63; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2114 = cache_hit ? _GEN_833 : valid_64; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2115 = cache_hit ? _GEN_834 : valid_65; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2116 = cache_hit ? _GEN_835 : valid_66; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2117 = cache_hit ? _GEN_836 : valid_67; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2118 = cache_hit ? _GEN_837 : valid_68; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2119 = cache_hit ? _GEN_838 : valid_69; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2120 = cache_hit ? _GEN_839 : valid_70; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2121 = cache_hit ? _GEN_840 : valid_71; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2122 = cache_hit ? _GEN_841 : valid_72; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2123 = cache_hit ? _GEN_842 : valid_73; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2124 = cache_hit ? _GEN_843 : valid_74; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2125 = cache_hit ? _GEN_844 : valid_75; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2126 = cache_hit ? _GEN_845 : valid_76; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2127 = cache_hit ? _GEN_846 : valid_77; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2128 = cache_hit ? _GEN_847 : valid_78; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2129 = cache_hit ? _GEN_848 : valid_79; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2130 = cache_hit ? _GEN_849 : valid_80; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2131 = cache_hit ? _GEN_850 : valid_81; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2132 = cache_hit ? _GEN_851 : valid_82; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2133 = cache_hit ? _GEN_852 : valid_83; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2134 = cache_hit ? _GEN_853 : valid_84; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2135 = cache_hit ? _GEN_854 : valid_85; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2136 = cache_hit ? _GEN_855 : valid_86; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2137 = cache_hit ? _GEN_856 : valid_87; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2138 = cache_hit ? _GEN_857 : valid_88; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2139 = cache_hit ? _GEN_858 : valid_89; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2140 = cache_hit ? _GEN_859 : valid_90; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2141 = cache_hit ? _GEN_860 : valid_91; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2142 = cache_hit ? _GEN_861 : valid_92; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2143 = cache_hit ? _GEN_862 : valid_93; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2144 = cache_hit ? _GEN_863 : valid_94; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2145 = cache_hit ? _GEN_864 : valid_95; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2146 = cache_hit ? _GEN_865 : valid_96; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2147 = cache_hit ? _GEN_866 : valid_97; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2148 = cache_hit ? _GEN_867 : valid_98; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2149 = cache_hit ? _GEN_868 : valid_99; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2150 = cache_hit ? _GEN_869 : valid_100; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2151 = cache_hit ? _GEN_870 : valid_101; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2152 = cache_hit ? _GEN_871 : valid_102; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2153 = cache_hit ? _GEN_872 : valid_103; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2154 = cache_hit ? _GEN_873 : valid_104; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2155 = cache_hit ? _GEN_874 : valid_105; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2156 = cache_hit ? _GEN_875 : valid_106; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2157 = cache_hit ? _GEN_876 : valid_107; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2158 = cache_hit ? _GEN_877 : valid_108; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2159 = cache_hit ? _GEN_878 : valid_109; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2160 = cache_hit ? _GEN_879 : valid_110; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2161 = cache_hit ? _GEN_880 : valid_111; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2162 = cache_hit ? _GEN_881 : valid_112; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2163 = cache_hit ? _GEN_882 : valid_113; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2164 = cache_hit ? _GEN_883 : valid_114; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2165 = cache_hit ? _GEN_884 : valid_115; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2166 = cache_hit ? _GEN_885 : valid_116; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2167 = cache_hit ? _GEN_886 : valid_117; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2168 = cache_hit ? _GEN_887 : valid_118; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2169 = cache_hit ? _GEN_888 : valid_119; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2170 = cache_hit ? _GEN_889 : valid_120; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2171 = cache_hit ? _GEN_890 : valid_121; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2172 = cache_hit ? _GEN_891 : valid_122; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2173 = cache_hit ? _GEN_892 : valid_123; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2174 = cache_hit ? _GEN_893 : valid_124; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2175 = cache_hit ? _GEN_894 : valid_125; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2176 = cache_hit ? _GEN_895 : valid_126; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2177 = cache_hit ? _GEN_896 : valid_127; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2178 = cache_hit ? _GEN_897 : valid_128; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2179 = cache_hit ? _GEN_898 : valid_129; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2180 = cache_hit ? _GEN_899 : valid_130; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2181 = cache_hit ? _GEN_900 : valid_131; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2182 = cache_hit ? _GEN_901 : valid_132; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2183 = cache_hit ? _GEN_902 : valid_133; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2184 = cache_hit ? _GEN_903 : valid_134; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2185 = cache_hit ? _GEN_904 : valid_135; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2186 = cache_hit ? _GEN_905 : valid_136; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2187 = cache_hit ? _GEN_906 : valid_137; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2188 = cache_hit ? _GEN_907 : valid_138; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2189 = cache_hit ? _GEN_908 : valid_139; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2190 = cache_hit ? _GEN_909 : valid_140; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2191 = cache_hit ? _GEN_910 : valid_141; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2192 = cache_hit ? _GEN_911 : valid_142; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2193 = cache_hit ? _GEN_912 : valid_143; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2194 = cache_hit ? _GEN_913 : valid_144; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2195 = cache_hit ? _GEN_914 : valid_145; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2196 = cache_hit ? _GEN_915 : valid_146; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2197 = cache_hit ? _GEN_916 : valid_147; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2198 = cache_hit ? _GEN_917 : valid_148; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2199 = cache_hit ? _GEN_918 : valid_149; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2200 = cache_hit ? _GEN_919 : valid_150; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2201 = cache_hit ? _GEN_920 : valid_151; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2202 = cache_hit ? _GEN_921 : valid_152; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2203 = cache_hit ? _GEN_922 : valid_153; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2204 = cache_hit ? _GEN_923 : valid_154; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2205 = cache_hit ? _GEN_924 : valid_155; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2206 = cache_hit ? _GEN_925 : valid_156; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2207 = cache_hit ? _GEN_926 : valid_157; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2208 = cache_hit ? _GEN_927 : valid_158; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2209 = cache_hit ? _GEN_928 : valid_159; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2210 = cache_hit ? _GEN_929 : valid_160; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2211 = cache_hit ? _GEN_930 : valid_161; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2212 = cache_hit ? _GEN_931 : valid_162; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2213 = cache_hit ? _GEN_932 : valid_163; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2214 = cache_hit ? _GEN_933 : valid_164; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2215 = cache_hit ? _GEN_934 : valid_165; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2216 = cache_hit ? _GEN_935 : valid_166; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2217 = cache_hit ? _GEN_936 : valid_167; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2218 = cache_hit ? _GEN_937 : valid_168; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2219 = cache_hit ? _GEN_938 : valid_169; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2220 = cache_hit ? _GEN_939 : valid_170; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2221 = cache_hit ? _GEN_940 : valid_171; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2222 = cache_hit ? _GEN_941 : valid_172; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2223 = cache_hit ? _GEN_942 : valid_173; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2224 = cache_hit ? _GEN_943 : valid_174; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2225 = cache_hit ? _GEN_944 : valid_175; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2226 = cache_hit ? _GEN_945 : valid_176; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2227 = cache_hit ? _GEN_946 : valid_177; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2228 = cache_hit ? _GEN_947 : valid_178; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2229 = cache_hit ? _GEN_948 : valid_179; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2230 = cache_hit ? _GEN_949 : valid_180; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2231 = cache_hit ? _GEN_950 : valid_181; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2232 = cache_hit ? _GEN_951 : valid_182; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2233 = cache_hit ? _GEN_952 : valid_183; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2234 = cache_hit ? _GEN_953 : valid_184; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2235 = cache_hit ? _GEN_954 : valid_185; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2236 = cache_hit ? _GEN_955 : valid_186; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2237 = cache_hit ? _GEN_956 : valid_187; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2238 = cache_hit ? _GEN_957 : valid_188; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2239 = cache_hit ? _GEN_958 : valid_189; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2240 = cache_hit ? _GEN_959 : valid_190; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2241 = cache_hit ? _GEN_960 : valid_191; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2242 = cache_hit ? _GEN_961 : valid_192; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2243 = cache_hit ? _GEN_962 : valid_193; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2244 = cache_hit ? _GEN_963 : valid_194; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2245 = cache_hit ? _GEN_964 : valid_195; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2246 = cache_hit ? _GEN_965 : valid_196; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2247 = cache_hit ? _GEN_966 : valid_197; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2248 = cache_hit ? _GEN_967 : valid_198; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2249 = cache_hit ? _GEN_968 : valid_199; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2250 = cache_hit ? _GEN_969 : valid_200; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2251 = cache_hit ? _GEN_970 : valid_201; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2252 = cache_hit ? _GEN_971 : valid_202; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2253 = cache_hit ? _GEN_972 : valid_203; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2254 = cache_hit ? _GEN_973 : valid_204; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2255 = cache_hit ? _GEN_974 : valid_205; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2256 = cache_hit ? _GEN_975 : valid_206; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2257 = cache_hit ? _GEN_976 : valid_207; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2258 = cache_hit ? _GEN_977 : valid_208; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2259 = cache_hit ? _GEN_978 : valid_209; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2260 = cache_hit ? _GEN_979 : valid_210; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2261 = cache_hit ? _GEN_980 : valid_211; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2262 = cache_hit ? _GEN_981 : valid_212; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2263 = cache_hit ? _GEN_982 : valid_213; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2264 = cache_hit ? _GEN_983 : valid_214; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2265 = cache_hit ? _GEN_984 : valid_215; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2266 = cache_hit ? _GEN_985 : valid_216; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2267 = cache_hit ? _GEN_986 : valid_217; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2268 = cache_hit ? _GEN_987 : valid_218; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2269 = cache_hit ? _GEN_988 : valid_219; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2270 = cache_hit ? _GEN_989 : valid_220; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2271 = cache_hit ? _GEN_990 : valid_221; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2272 = cache_hit ? _GEN_991 : valid_222; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2273 = cache_hit ? _GEN_992 : valid_223; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2274 = cache_hit ? _GEN_993 : valid_224; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2275 = cache_hit ? _GEN_994 : valid_225; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2276 = cache_hit ? _GEN_995 : valid_226; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2277 = cache_hit ? _GEN_996 : valid_227; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2278 = cache_hit ? _GEN_997 : valid_228; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2279 = cache_hit ? _GEN_998 : valid_229; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2280 = cache_hit ? _GEN_999 : valid_230; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2281 = cache_hit ? _GEN_1000 : valid_231; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2282 = cache_hit ? _GEN_1001 : valid_232; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2283 = cache_hit ? _GEN_1002 : valid_233; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2284 = cache_hit ? _GEN_1003 : valid_234; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2285 = cache_hit ? _GEN_1004 : valid_235; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2286 = cache_hit ? _GEN_1005 : valid_236; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2287 = cache_hit ? _GEN_1006 : valid_237; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2288 = cache_hit ? _GEN_1007 : valid_238; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2289 = cache_hit ? _GEN_1008 : valid_239; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2290 = cache_hit ? _GEN_1009 : valid_240; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2291 = cache_hit ? _GEN_1010 : valid_241; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2292 = cache_hit ? _GEN_1011 : valid_242; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2293 = cache_hit ? _GEN_1012 : valid_243; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2294 = cache_hit ? _GEN_1013 : valid_244; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2295 = cache_hit ? _GEN_1014 : valid_245; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2296 = cache_hit ? _GEN_1015 : valid_246; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2297 = cache_hit ? _GEN_1016 : valid_247; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2298 = cache_hit ? _GEN_1017 : valid_248; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2299 = cache_hit ? _GEN_1018 : valid_249; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2300 = cache_hit ? _GEN_1019 : valid_250; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2301 = cache_hit ? _GEN_1020 : valid_251; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2302 = cache_hit ? _GEN_1021 : valid_252; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2303 = cache_hit ? _GEN_1022 : valid_253; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2304 = cache_hit ? _GEN_1023 : valid_254; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire  _GEN_2305 = cache_hit ? _GEN_1024 : valid_255; // @[Dcache.scala 134:29 Dcache.scala 17:24]
  wire [19:0] _GEN_2306 = cache_hit ? _GEN_1025 : tag_0; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2307 = cache_hit ? _GEN_1026 : tag_1; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2308 = cache_hit ? _GEN_1027 : tag_2; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2309 = cache_hit ? _GEN_1028 : tag_3; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2310 = cache_hit ? _GEN_1029 : tag_4; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2311 = cache_hit ? _GEN_1030 : tag_5; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2312 = cache_hit ? _GEN_1031 : tag_6; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2313 = cache_hit ? _GEN_1032 : tag_7; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2314 = cache_hit ? _GEN_1033 : tag_8; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2315 = cache_hit ? _GEN_1034 : tag_9; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2316 = cache_hit ? _GEN_1035 : tag_10; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2317 = cache_hit ? _GEN_1036 : tag_11; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2318 = cache_hit ? _GEN_1037 : tag_12; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2319 = cache_hit ? _GEN_1038 : tag_13; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2320 = cache_hit ? _GEN_1039 : tag_14; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2321 = cache_hit ? _GEN_1040 : tag_15; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2322 = cache_hit ? _GEN_1041 : tag_16; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2323 = cache_hit ? _GEN_1042 : tag_17; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2324 = cache_hit ? _GEN_1043 : tag_18; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2325 = cache_hit ? _GEN_1044 : tag_19; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2326 = cache_hit ? _GEN_1045 : tag_20; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2327 = cache_hit ? _GEN_1046 : tag_21; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2328 = cache_hit ? _GEN_1047 : tag_22; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2329 = cache_hit ? _GEN_1048 : tag_23; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2330 = cache_hit ? _GEN_1049 : tag_24; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2331 = cache_hit ? _GEN_1050 : tag_25; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2332 = cache_hit ? _GEN_1051 : tag_26; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2333 = cache_hit ? _GEN_1052 : tag_27; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2334 = cache_hit ? _GEN_1053 : tag_28; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2335 = cache_hit ? _GEN_1054 : tag_29; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2336 = cache_hit ? _GEN_1055 : tag_30; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2337 = cache_hit ? _GEN_1056 : tag_31; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2338 = cache_hit ? _GEN_1057 : tag_32; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2339 = cache_hit ? _GEN_1058 : tag_33; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2340 = cache_hit ? _GEN_1059 : tag_34; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2341 = cache_hit ? _GEN_1060 : tag_35; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2342 = cache_hit ? _GEN_1061 : tag_36; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2343 = cache_hit ? _GEN_1062 : tag_37; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2344 = cache_hit ? _GEN_1063 : tag_38; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2345 = cache_hit ? _GEN_1064 : tag_39; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2346 = cache_hit ? _GEN_1065 : tag_40; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2347 = cache_hit ? _GEN_1066 : tag_41; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2348 = cache_hit ? _GEN_1067 : tag_42; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2349 = cache_hit ? _GEN_1068 : tag_43; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2350 = cache_hit ? _GEN_1069 : tag_44; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2351 = cache_hit ? _GEN_1070 : tag_45; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2352 = cache_hit ? _GEN_1071 : tag_46; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2353 = cache_hit ? _GEN_1072 : tag_47; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2354 = cache_hit ? _GEN_1073 : tag_48; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2355 = cache_hit ? _GEN_1074 : tag_49; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2356 = cache_hit ? _GEN_1075 : tag_50; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2357 = cache_hit ? _GEN_1076 : tag_51; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2358 = cache_hit ? _GEN_1077 : tag_52; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2359 = cache_hit ? _GEN_1078 : tag_53; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2360 = cache_hit ? _GEN_1079 : tag_54; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2361 = cache_hit ? _GEN_1080 : tag_55; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2362 = cache_hit ? _GEN_1081 : tag_56; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2363 = cache_hit ? _GEN_1082 : tag_57; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2364 = cache_hit ? _GEN_1083 : tag_58; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2365 = cache_hit ? _GEN_1084 : tag_59; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2366 = cache_hit ? _GEN_1085 : tag_60; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2367 = cache_hit ? _GEN_1086 : tag_61; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2368 = cache_hit ? _GEN_1087 : tag_62; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2369 = cache_hit ? _GEN_1088 : tag_63; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2370 = cache_hit ? _GEN_1089 : tag_64; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2371 = cache_hit ? _GEN_1090 : tag_65; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2372 = cache_hit ? _GEN_1091 : tag_66; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2373 = cache_hit ? _GEN_1092 : tag_67; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2374 = cache_hit ? _GEN_1093 : tag_68; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2375 = cache_hit ? _GEN_1094 : tag_69; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2376 = cache_hit ? _GEN_1095 : tag_70; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2377 = cache_hit ? _GEN_1096 : tag_71; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2378 = cache_hit ? _GEN_1097 : tag_72; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2379 = cache_hit ? _GEN_1098 : tag_73; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2380 = cache_hit ? _GEN_1099 : tag_74; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2381 = cache_hit ? _GEN_1100 : tag_75; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2382 = cache_hit ? _GEN_1101 : tag_76; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2383 = cache_hit ? _GEN_1102 : tag_77; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2384 = cache_hit ? _GEN_1103 : tag_78; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2385 = cache_hit ? _GEN_1104 : tag_79; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2386 = cache_hit ? _GEN_1105 : tag_80; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2387 = cache_hit ? _GEN_1106 : tag_81; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2388 = cache_hit ? _GEN_1107 : tag_82; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2389 = cache_hit ? _GEN_1108 : tag_83; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2390 = cache_hit ? _GEN_1109 : tag_84; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2391 = cache_hit ? _GEN_1110 : tag_85; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2392 = cache_hit ? _GEN_1111 : tag_86; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2393 = cache_hit ? _GEN_1112 : tag_87; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2394 = cache_hit ? _GEN_1113 : tag_88; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2395 = cache_hit ? _GEN_1114 : tag_89; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2396 = cache_hit ? _GEN_1115 : tag_90; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2397 = cache_hit ? _GEN_1116 : tag_91; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2398 = cache_hit ? _GEN_1117 : tag_92; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2399 = cache_hit ? _GEN_1118 : tag_93; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2400 = cache_hit ? _GEN_1119 : tag_94; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2401 = cache_hit ? _GEN_1120 : tag_95; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2402 = cache_hit ? _GEN_1121 : tag_96; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2403 = cache_hit ? _GEN_1122 : tag_97; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2404 = cache_hit ? _GEN_1123 : tag_98; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2405 = cache_hit ? _GEN_1124 : tag_99; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2406 = cache_hit ? _GEN_1125 : tag_100; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2407 = cache_hit ? _GEN_1126 : tag_101; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2408 = cache_hit ? _GEN_1127 : tag_102; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2409 = cache_hit ? _GEN_1128 : tag_103; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2410 = cache_hit ? _GEN_1129 : tag_104; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2411 = cache_hit ? _GEN_1130 : tag_105; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2412 = cache_hit ? _GEN_1131 : tag_106; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2413 = cache_hit ? _GEN_1132 : tag_107; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2414 = cache_hit ? _GEN_1133 : tag_108; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2415 = cache_hit ? _GEN_1134 : tag_109; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2416 = cache_hit ? _GEN_1135 : tag_110; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2417 = cache_hit ? _GEN_1136 : tag_111; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2418 = cache_hit ? _GEN_1137 : tag_112; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2419 = cache_hit ? _GEN_1138 : tag_113; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2420 = cache_hit ? _GEN_1139 : tag_114; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2421 = cache_hit ? _GEN_1140 : tag_115; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2422 = cache_hit ? _GEN_1141 : tag_116; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2423 = cache_hit ? _GEN_1142 : tag_117; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2424 = cache_hit ? _GEN_1143 : tag_118; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2425 = cache_hit ? _GEN_1144 : tag_119; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2426 = cache_hit ? _GEN_1145 : tag_120; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2427 = cache_hit ? _GEN_1146 : tag_121; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2428 = cache_hit ? _GEN_1147 : tag_122; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2429 = cache_hit ? _GEN_1148 : tag_123; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2430 = cache_hit ? _GEN_1149 : tag_124; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2431 = cache_hit ? _GEN_1150 : tag_125; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2432 = cache_hit ? _GEN_1151 : tag_126; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2433 = cache_hit ? _GEN_1152 : tag_127; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2434 = cache_hit ? _GEN_1153 : tag_128; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2435 = cache_hit ? _GEN_1154 : tag_129; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2436 = cache_hit ? _GEN_1155 : tag_130; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2437 = cache_hit ? _GEN_1156 : tag_131; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2438 = cache_hit ? _GEN_1157 : tag_132; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2439 = cache_hit ? _GEN_1158 : tag_133; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2440 = cache_hit ? _GEN_1159 : tag_134; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2441 = cache_hit ? _GEN_1160 : tag_135; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2442 = cache_hit ? _GEN_1161 : tag_136; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2443 = cache_hit ? _GEN_1162 : tag_137; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2444 = cache_hit ? _GEN_1163 : tag_138; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2445 = cache_hit ? _GEN_1164 : tag_139; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2446 = cache_hit ? _GEN_1165 : tag_140; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2447 = cache_hit ? _GEN_1166 : tag_141; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2448 = cache_hit ? _GEN_1167 : tag_142; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2449 = cache_hit ? _GEN_1168 : tag_143; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2450 = cache_hit ? _GEN_1169 : tag_144; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2451 = cache_hit ? _GEN_1170 : tag_145; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2452 = cache_hit ? _GEN_1171 : tag_146; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2453 = cache_hit ? _GEN_1172 : tag_147; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2454 = cache_hit ? _GEN_1173 : tag_148; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2455 = cache_hit ? _GEN_1174 : tag_149; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2456 = cache_hit ? _GEN_1175 : tag_150; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2457 = cache_hit ? _GEN_1176 : tag_151; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2458 = cache_hit ? _GEN_1177 : tag_152; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2459 = cache_hit ? _GEN_1178 : tag_153; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2460 = cache_hit ? _GEN_1179 : tag_154; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2461 = cache_hit ? _GEN_1180 : tag_155; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2462 = cache_hit ? _GEN_1181 : tag_156; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2463 = cache_hit ? _GEN_1182 : tag_157; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2464 = cache_hit ? _GEN_1183 : tag_158; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2465 = cache_hit ? _GEN_1184 : tag_159; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2466 = cache_hit ? _GEN_1185 : tag_160; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2467 = cache_hit ? _GEN_1186 : tag_161; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2468 = cache_hit ? _GEN_1187 : tag_162; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2469 = cache_hit ? _GEN_1188 : tag_163; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2470 = cache_hit ? _GEN_1189 : tag_164; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2471 = cache_hit ? _GEN_1190 : tag_165; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2472 = cache_hit ? _GEN_1191 : tag_166; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2473 = cache_hit ? _GEN_1192 : tag_167; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2474 = cache_hit ? _GEN_1193 : tag_168; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2475 = cache_hit ? _GEN_1194 : tag_169; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2476 = cache_hit ? _GEN_1195 : tag_170; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2477 = cache_hit ? _GEN_1196 : tag_171; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2478 = cache_hit ? _GEN_1197 : tag_172; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2479 = cache_hit ? _GEN_1198 : tag_173; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2480 = cache_hit ? _GEN_1199 : tag_174; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2481 = cache_hit ? _GEN_1200 : tag_175; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2482 = cache_hit ? _GEN_1201 : tag_176; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2483 = cache_hit ? _GEN_1202 : tag_177; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2484 = cache_hit ? _GEN_1203 : tag_178; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2485 = cache_hit ? _GEN_1204 : tag_179; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2486 = cache_hit ? _GEN_1205 : tag_180; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2487 = cache_hit ? _GEN_1206 : tag_181; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2488 = cache_hit ? _GEN_1207 : tag_182; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2489 = cache_hit ? _GEN_1208 : tag_183; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2490 = cache_hit ? _GEN_1209 : tag_184; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2491 = cache_hit ? _GEN_1210 : tag_185; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2492 = cache_hit ? _GEN_1211 : tag_186; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2493 = cache_hit ? _GEN_1212 : tag_187; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2494 = cache_hit ? _GEN_1213 : tag_188; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2495 = cache_hit ? _GEN_1214 : tag_189; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2496 = cache_hit ? _GEN_1215 : tag_190; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2497 = cache_hit ? _GEN_1216 : tag_191; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2498 = cache_hit ? _GEN_1217 : tag_192; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2499 = cache_hit ? _GEN_1218 : tag_193; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2500 = cache_hit ? _GEN_1219 : tag_194; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2501 = cache_hit ? _GEN_1220 : tag_195; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2502 = cache_hit ? _GEN_1221 : tag_196; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2503 = cache_hit ? _GEN_1222 : tag_197; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2504 = cache_hit ? _GEN_1223 : tag_198; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2505 = cache_hit ? _GEN_1224 : tag_199; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2506 = cache_hit ? _GEN_1225 : tag_200; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2507 = cache_hit ? _GEN_1226 : tag_201; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2508 = cache_hit ? _GEN_1227 : tag_202; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2509 = cache_hit ? _GEN_1228 : tag_203; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2510 = cache_hit ? _GEN_1229 : tag_204; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2511 = cache_hit ? _GEN_1230 : tag_205; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2512 = cache_hit ? _GEN_1231 : tag_206; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2513 = cache_hit ? _GEN_1232 : tag_207; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2514 = cache_hit ? _GEN_1233 : tag_208; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2515 = cache_hit ? _GEN_1234 : tag_209; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2516 = cache_hit ? _GEN_1235 : tag_210; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2517 = cache_hit ? _GEN_1236 : tag_211; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2518 = cache_hit ? _GEN_1237 : tag_212; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2519 = cache_hit ? _GEN_1238 : tag_213; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2520 = cache_hit ? _GEN_1239 : tag_214; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2521 = cache_hit ? _GEN_1240 : tag_215; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2522 = cache_hit ? _GEN_1241 : tag_216; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2523 = cache_hit ? _GEN_1242 : tag_217; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2524 = cache_hit ? _GEN_1243 : tag_218; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2525 = cache_hit ? _GEN_1244 : tag_219; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2526 = cache_hit ? _GEN_1245 : tag_220; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2527 = cache_hit ? _GEN_1246 : tag_221; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2528 = cache_hit ? _GEN_1247 : tag_222; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2529 = cache_hit ? _GEN_1248 : tag_223; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2530 = cache_hit ? _GEN_1249 : tag_224; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2531 = cache_hit ? _GEN_1250 : tag_225; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2532 = cache_hit ? _GEN_1251 : tag_226; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2533 = cache_hit ? _GEN_1252 : tag_227; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2534 = cache_hit ? _GEN_1253 : tag_228; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2535 = cache_hit ? _GEN_1254 : tag_229; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2536 = cache_hit ? _GEN_1255 : tag_230; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2537 = cache_hit ? _GEN_1256 : tag_231; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2538 = cache_hit ? _GEN_1257 : tag_232; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2539 = cache_hit ? _GEN_1258 : tag_233; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2540 = cache_hit ? _GEN_1259 : tag_234; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2541 = cache_hit ? _GEN_1260 : tag_235; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2542 = cache_hit ? _GEN_1261 : tag_236; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2543 = cache_hit ? _GEN_1262 : tag_237; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2544 = cache_hit ? _GEN_1263 : tag_238; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2545 = cache_hit ? _GEN_1264 : tag_239; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2546 = cache_hit ? _GEN_1265 : tag_240; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2547 = cache_hit ? _GEN_1266 : tag_241; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2548 = cache_hit ? _GEN_1267 : tag_242; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2549 = cache_hit ? _GEN_1268 : tag_243; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2550 = cache_hit ? _GEN_1269 : tag_244; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2551 = cache_hit ? _GEN_1270 : tag_245; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2552 = cache_hit ? _GEN_1271 : tag_246; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2553 = cache_hit ? _GEN_1272 : tag_247; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2554 = cache_hit ? _GEN_1273 : tag_248; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2555 = cache_hit ? _GEN_1274 : tag_249; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2556 = cache_hit ? _GEN_1275 : tag_250; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2557 = cache_hit ? _GEN_1276 : tag_251; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2558 = cache_hit ? _GEN_1277 : tag_252; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2559 = cache_hit ? _GEN_1278 : tag_253; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2560 = cache_hit ? _GEN_1279 : tag_254; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [19:0] _GEN_2561 = cache_hit ? _GEN_1280 : tag_255; // @[Dcache.scala 134:29 Dcache.scala 16:24]
  wire [3:0] _GEN_2562 = cache_hit ? _GEN_1281 : offset_0; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2563 = cache_hit ? _GEN_1282 : offset_1; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2564 = cache_hit ? _GEN_1283 : offset_2; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2565 = cache_hit ? _GEN_1284 : offset_3; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2566 = cache_hit ? _GEN_1285 : offset_4; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2567 = cache_hit ? _GEN_1286 : offset_5; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2568 = cache_hit ? _GEN_1287 : offset_6; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2569 = cache_hit ? _GEN_1288 : offset_7; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2570 = cache_hit ? _GEN_1289 : offset_8; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2571 = cache_hit ? _GEN_1290 : offset_9; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2572 = cache_hit ? _GEN_1291 : offset_10; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2573 = cache_hit ? _GEN_1292 : offset_11; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2574 = cache_hit ? _GEN_1293 : offset_12; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2575 = cache_hit ? _GEN_1294 : offset_13; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2576 = cache_hit ? _GEN_1295 : offset_14; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2577 = cache_hit ? _GEN_1296 : offset_15; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2578 = cache_hit ? _GEN_1297 : offset_16; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2579 = cache_hit ? _GEN_1298 : offset_17; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2580 = cache_hit ? _GEN_1299 : offset_18; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2581 = cache_hit ? _GEN_1300 : offset_19; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2582 = cache_hit ? _GEN_1301 : offset_20; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2583 = cache_hit ? _GEN_1302 : offset_21; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2584 = cache_hit ? _GEN_1303 : offset_22; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2585 = cache_hit ? _GEN_1304 : offset_23; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2586 = cache_hit ? _GEN_1305 : offset_24; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2587 = cache_hit ? _GEN_1306 : offset_25; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2588 = cache_hit ? _GEN_1307 : offset_26; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2589 = cache_hit ? _GEN_1308 : offset_27; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2590 = cache_hit ? _GEN_1309 : offset_28; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2591 = cache_hit ? _GEN_1310 : offset_29; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2592 = cache_hit ? _GEN_1311 : offset_30; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2593 = cache_hit ? _GEN_1312 : offset_31; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2594 = cache_hit ? _GEN_1313 : offset_32; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2595 = cache_hit ? _GEN_1314 : offset_33; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2596 = cache_hit ? _GEN_1315 : offset_34; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2597 = cache_hit ? _GEN_1316 : offset_35; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2598 = cache_hit ? _GEN_1317 : offset_36; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2599 = cache_hit ? _GEN_1318 : offset_37; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2600 = cache_hit ? _GEN_1319 : offset_38; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2601 = cache_hit ? _GEN_1320 : offset_39; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2602 = cache_hit ? _GEN_1321 : offset_40; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2603 = cache_hit ? _GEN_1322 : offset_41; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2604 = cache_hit ? _GEN_1323 : offset_42; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2605 = cache_hit ? _GEN_1324 : offset_43; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2606 = cache_hit ? _GEN_1325 : offset_44; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2607 = cache_hit ? _GEN_1326 : offset_45; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2608 = cache_hit ? _GEN_1327 : offset_46; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2609 = cache_hit ? _GEN_1328 : offset_47; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2610 = cache_hit ? _GEN_1329 : offset_48; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2611 = cache_hit ? _GEN_1330 : offset_49; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2612 = cache_hit ? _GEN_1331 : offset_50; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2613 = cache_hit ? _GEN_1332 : offset_51; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2614 = cache_hit ? _GEN_1333 : offset_52; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2615 = cache_hit ? _GEN_1334 : offset_53; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2616 = cache_hit ? _GEN_1335 : offset_54; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2617 = cache_hit ? _GEN_1336 : offset_55; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2618 = cache_hit ? _GEN_1337 : offset_56; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2619 = cache_hit ? _GEN_1338 : offset_57; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2620 = cache_hit ? _GEN_1339 : offset_58; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2621 = cache_hit ? _GEN_1340 : offset_59; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2622 = cache_hit ? _GEN_1341 : offset_60; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2623 = cache_hit ? _GEN_1342 : offset_61; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2624 = cache_hit ? _GEN_1343 : offset_62; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2625 = cache_hit ? _GEN_1344 : offset_63; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2626 = cache_hit ? _GEN_1345 : offset_64; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2627 = cache_hit ? _GEN_1346 : offset_65; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2628 = cache_hit ? _GEN_1347 : offset_66; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2629 = cache_hit ? _GEN_1348 : offset_67; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2630 = cache_hit ? _GEN_1349 : offset_68; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2631 = cache_hit ? _GEN_1350 : offset_69; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2632 = cache_hit ? _GEN_1351 : offset_70; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2633 = cache_hit ? _GEN_1352 : offset_71; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2634 = cache_hit ? _GEN_1353 : offset_72; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2635 = cache_hit ? _GEN_1354 : offset_73; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2636 = cache_hit ? _GEN_1355 : offset_74; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2637 = cache_hit ? _GEN_1356 : offset_75; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2638 = cache_hit ? _GEN_1357 : offset_76; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2639 = cache_hit ? _GEN_1358 : offset_77; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2640 = cache_hit ? _GEN_1359 : offset_78; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2641 = cache_hit ? _GEN_1360 : offset_79; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2642 = cache_hit ? _GEN_1361 : offset_80; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2643 = cache_hit ? _GEN_1362 : offset_81; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2644 = cache_hit ? _GEN_1363 : offset_82; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2645 = cache_hit ? _GEN_1364 : offset_83; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2646 = cache_hit ? _GEN_1365 : offset_84; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2647 = cache_hit ? _GEN_1366 : offset_85; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2648 = cache_hit ? _GEN_1367 : offset_86; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2649 = cache_hit ? _GEN_1368 : offset_87; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2650 = cache_hit ? _GEN_1369 : offset_88; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2651 = cache_hit ? _GEN_1370 : offset_89; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2652 = cache_hit ? _GEN_1371 : offset_90; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2653 = cache_hit ? _GEN_1372 : offset_91; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2654 = cache_hit ? _GEN_1373 : offset_92; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2655 = cache_hit ? _GEN_1374 : offset_93; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2656 = cache_hit ? _GEN_1375 : offset_94; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2657 = cache_hit ? _GEN_1376 : offset_95; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2658 = cache_hit ? _GEN_1377 : offset_96; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2659 = cache_hit ? _GEN_1378 : offset_97; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2660 = cache_hit ? _GEN_1379 : offset_98; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2661 = cache_hit ? _GEN_1380 : offset_99; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2662 = cache_hit ? _GEN_1381 : offset_100; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2663 = cache_hit ? _GEN_1382 : offset_101; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2664 = cache_hit ? _GEN_1383 : offset_102; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2665 = cache_hit ? _GEN_1384 : offset_103; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2666 = cache_hit ? _GEN_1385 : offset_104; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2667 = cache_hit ? _GEN_1386 : offset_105; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2668 = cache_hit ? _GEN_1387 : offset_106; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2669 = cache_hit ? _GEN_1388 : offset_107; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2670 = cache_hit ? _GEN_1389 : offset_108; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2671 = cache_hit ? _GEN_1390 : offset_109; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2672 = cache_hit ? _GEN_1391 : offset_110; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2673 = cache_hit ? _GEN_1392 : offset_111; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2674 = cache_hit ? _GEN_1393 : offset_112; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2675 = cache_hit ? _GEN_1394 : offset_113; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2676 = cache_hit ? _GEN_1395 : offset_114; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2677 = cache_hit ? _GEN_1396 : offset_115; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2678 = cache_hit ? _GEN_1397 : offset_116; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2679 = cache_hit ? _GEN_1398 : offset_117; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2680 = cache_hit ? _GEN_1399 : offset_118; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2681 = cache_hit ? _GEN_1400 : offset_119; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2682 = cache_hit ? _GEN_1401 : offset_120; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2683 = cache_hit ? _GEN_1402 : offset_121; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2684 = cache_hit ? _GEN_1403 : offset_122; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2685 = cache_hit ? _GEN_1404 : offset_123; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2686 = cache_hit ? _GEN_1405 : offset_124; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2687 = cache_hit ? _GEN_1406 : offset_125; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2688 = cache_hit ? _GEN_1407 : offset_126; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2689 = cache_hit ? _GEN_1408 : offset_127; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2690 = cache_hit ? _GEN_1409 : offset_128; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2691 = cache_hit ? _GEN_1410 : offset_129; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2692 = cache_hit ? _GEN_1411 : offset_130; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2693 = cache_hit ? _GEN_1412 : offset_131; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2694 = cache_hit ? _GEN_1413 : offset_132; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2695 = cache_hit ? _GEN_1414 : offset_133; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2696 = cache_hit ? _GEN_1415 : offset_134; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2697 = cache_hit ? _GEN_1416 : offset_135; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2698 = cache_hit ? _GEN_1417 : offset_136; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2699 = cache_hit ? _GEN_1418 : offset_137; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2700 = cache_hit ? _GEN_1419 : offset_138; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2701 = cache_hit ? _GEN_1420 : offset_139; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2702 = cache_hit ? _GEN_1421 : offset_140; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2703 = cache_hit ? _GEN_1422 : offset_141; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2704 = cache_hit ? _GEN_1423 : offset_142; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2705 = cache_hit ? _GEN_1424 : offset_143; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2706 = cache_hit ? _GEN_1425 : offset_144; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2707 = cache_hit ? _GEN_1426 : offset_145; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2708 = cache_hit ? _GEN_1427 : offset_146; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2709 = cache_hit ? _GEN_1428 : offset_147; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2710 = cache_hit ? _GEN_1429 : offset_148; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2711 = cache_hit ? _GEN_1430 : offset_149; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2712 = cache_hit ? _GEN_1431 : offset_150; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2713 = cache_hit ? _GEN_1432 : offset_151; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2714 = cache_hit ? _GEN_1433 : offset_152; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2715 = cache_hit ? _GEN_1434 : offset_153; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2716 = cache_hit ? _GEN_1435 : offset_154; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2717 = cache_hit ? _GEN_1436 : offset_155; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2718 = cache_hit ? _GEN_1437 : offset_156; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2719 = cache_hit ? _GEN_1438 : offset_157; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2720 = cache_hit ? _GEN_1439 : offset_158; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2721 = cache_hit ? _GEN_1440 : offset_159; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2722 = cache_hit ? _GEN_1441 : offset_160; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2723 = cache_hit ? _GEN_1442 : offset_161; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2724 = cache_hit ? _GEN_1443 : offset_162; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2725 = cache_hit ? _GEN_1444 : offset_163; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2726 = cache_hit ? _GEN_1445 : offset_164; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2727 = cache_hit ? _GEN_1446 : offset_165; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2728 = cache_hit ? _GEN_1447 : offset_166; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2729 = cache_hit ? _GEN_1448 : offset_167; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2730 = cache_hit ? _GEN_1449 : offset_168; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2731 = cache_hit ? _GEN_1450 : offset_169; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2732 = cache_hit ? _GEN_1451 : offset_170; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2733 = cache_hit ? _GEN_1452 : offset_171; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2734 = cache_hit ? _GEN_1453 : offset_172; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2735 = cache_hit ? _GEN_1454 : offset_173; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2736 = cache_hit ? _GEN_1455 : offset_174; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2737 = cache_hit ? _GEN_1456 : offset_175; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2738 = cache_hit ? _GEN_1457 : offset_176; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2739 = cache_hit ? _GEN_1458 : offset_177; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2740 = cache_hit ? _GEN_1459 : offset_178; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2741 = cache_hit ? _GEN_1460 : offset_179; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2742 = cache_hit ? _GEN_1461 : offset_180; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2743 = cache_hit ? _GEN_1462 : offset_181; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2744 = cache_hit ? _GEN_1463 : offset_182; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2745 = cache_hit ? _GEN_1464 : offset_183; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2746 = cache_hit ? _GEN_1465 : offset_184; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2747 = cache_hit ? _GEN_1466 : offset_185; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2748 = cache_hit ? _GEN_1467 : offset_186; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2749 = cache_hit ? _GEN_1468 : offset_187; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2750 = cache_hit ? _GEN_1469 : offset_188; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2751 = cache_hit ? _GEN_1470 : offset_189; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2752 = cache_hit ? _GEN_1471 : offset_190; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2753 = cache_hit ? _GEN_1472 : offset_191; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2754 = cache_hit ? _GEN_1473 : offset_192; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2755 = cache_hit ? _GEN_1474 : offset_193; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2756 = cache_hit ? _GEN_1475 : offset_194; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2757 = cache_hit ? _GEN_1476 : offset_195; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2758 = cache_hit ? _GEN_1477 : offset_196; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2759 = cache_hit ? _GEN_1478 : offset_197; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2760 = cache_hit ? _GEN_1479 : offset_198; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2761 = cache_hit ? _GEN_1480 : offset_199; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2762 = cache_hit ? _GEN_1481 : offset_200; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2763 = cache_hit ? _GEN_1482 : offset_201; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2764 = cache_hit ? _GEN_1483 : offset_202; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2765 = cache_hit ? _GEN_1484 : offset_203; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2766 = cache_hit ? _GEN_1485 : offset_204; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2767 = cache_hit ? _GEN_1486 : offset_205; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2768 = cache_hit ? _GEN_1487 : offset_206; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2769 = cache_hit ? _GEN_1488 : offset_207; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2770 = cache_hit ? _GEN_1489 : offset_208; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2771 = cache_hit ? _GEN_1490 : offset_209; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2772 = cache_hit ? _GEN_1491 : offset_210; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2773 = cache_hit ? _GEN_1492 : offset_211; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2774 = cache_hit ? _GEN_1493 : offset_212; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2775 = cache_hit ? _GEN_1494 : offset_213; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2776 = cache_hit ? _GEN_1495 : offset_214; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2777 = cache_hit ? _GEN_1496 : offset_215; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2778 = cache_hit ? _GEN_1497 : offset_216; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2779 = cache_hit ? _GEN_1498 : offset_217; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2780 = cache_hit ? _GEN_1499 : offset_218; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2781 = cache_hit ? _GEN_1500 : offset_219; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2782 = cache_hit ? _GEN_1501 : offset_220; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2783 = cache_hit ? _GEN_1502 : offset_221; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2784 = cache_hit ? _GEN_1503 : offset_222; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2785 = cache_hit ? _GEN_1504 : offset_223; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2786 = cache_hit ? _GEN_1505 : offset_224; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2787 = cache_hit ? _GEN_1506 : offset_225; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2788 = cache_hit ? _GEN_1507 : offset_226; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2789 = cache_hit ? _GEN_1508 : offset_227; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2790 = cache_hit ? _GEN_1509 : offset_228; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2791 = cache_hit ? _GEN_1510 : offset_229; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2792 = cache_hit ? _GEN_1511 : offset_230; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2793 = cache_hit ? _GEN_1512 : offset_231; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2794 = cache_hit ? _GEN_1513 : offset_232; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2795 = cache_hit ? _GEN_1514 : offset_233; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2796 = cache_hit ? _GEN_1515 : offset_234; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2797 = cache_hit ? _GEN_1516 : offset_235; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2798 = cache_hit ? _GEN_1517 : offset_236; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2799 = cache_hit ? _GEN_1518 : offset_237; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2800 = cache_hit ? _GEN_1519 : offset_238; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2801 = cache_hit ? _GEN_1520 : offset_239; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2802 = cache_hit ? _GEN_1521 : offset_240; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2803 = cache_hit ? _GEN_1522 : offset_241; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2804 = cache_hit ? _GEN_1523 : offset_242; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2805 = cache_hit ? _GEN_1524 : offset_243; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2806 = cache_hit ? _GEN_1525 : offset_244; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2807 = cache_hit ? _GEN_1526 : offset_245; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2808 = cache_hit ? _GEN_1527 : offset_246; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2809 = cache_hit ? _GEN_1528 : offset_247; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2810 = cache_hit ? _GEN_1529 : offset_248; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2811 = cache_hit ? _GEN_1530 : offset_249; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2812 = cache_hit ? _GEN_1531 : offset_250; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2813 = cache_hit ? _GEN_1532 : offset_251; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2814 = cache_hit ? _GEN_1533 : offset_252; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2815 = cache_hit ? _GEN_1534 : offset_253; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2816 = cache_hit ? _GEN_1535 : offset_254; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire [3:0] _GEN_2817 = cache_hit ? _GEN_1536 : offset_255; // @[Dcache.scala 134:29 Dcache.scala 19:24]
  wire  _GEN_2818 = cache_hit | data_ready; // @[Dcache.scala 134:29 Dcache.scala 138:27 Dcache.scala 46:28]
  wire  _GEN_2819 = cache_hit ? io_dmem_data_req : cache_wen; // @[Dcache.scala 134:29 Dcache.scala 139:27 Dcache.scala 117:28]
  wire [127:0] _GEN_2820 = cache_hit ? _cache_wdata_T_3 : cache_wdata; // @[Dcache.scala 134:29 Dcache.scala 140:27 Dcache.scala 118:28]
  wire [127:0] _GEN_2821 = cache_hit ? _cache_strb_T_3 : cache_strb; // @[Dcache.scala 134:29 Dcache.scala 141:27 Dcache.scala 119:28]
  wire  _GEN_2822 = cache_hit ? _GEN_1793 : dirty_0; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2823 = cache_hit ? _GEN_1794 : dirty_1; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2824 = cache_hit ? _GEN_1795 : dirty_2; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2825 = cache_hit ? _GEN_1796 : dirty_3; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2826 = cache_hit ? _GEN_1797 : dirty_4; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2827 = cache_hit ? _GEN_1798 : dirty_5; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2828 = cache_hit ? _GEN_1799 : dirty_6; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2829 = cache_hit ? _GEN_1800 : dirty_7; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2830 = cache_hit ? _GEN_1801 : dirty_8; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2831 = cache_hit ? _GEN_1802 : dirty_9; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2832 = cache_hit ? _GEN_1803 : dirty_10; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2833 = cache_hit ? _GEN_1804 : dirty_11; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2834 = cache_hit ? _GEN_1805 : dirty_12; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2835 = cache_hit ? _GEN_1806 : dirty_13; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2836 = cache_hit ? _GEN_1807 : dirty_14; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2837 = cache_hit ? _GEN_1808 : dirty_15; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2838 = cache_hit ? _GEN_1809 : dirty_16; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2839 = cache_hit ? _GEN_1810 : dirty_17; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2840 = cache_hit ? _GEN_1811 : dirty_18; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2841 = cache_hit ? _GEN_1812 : dirty_19; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2842 = cache_hit ? _GEN_1813 : dirty_20; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2843 = cache_hit ? _GEN_1814 : dirty_21; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2844 = cache_hit ? _GEN_1815 : dirty_22; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2845 = cache_hit ? _GEN_1816 : dirty_23; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2846 = cache_hit ? _GEN_1817 : dirty_24; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2847 = cache_hit ? _GEN_1818 : dirty_25; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2848 = cache_hit ? _GEN_1819 : dirty_26; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2849 = cache_hit ? _GEN_1820 : dirty_27; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2850 = cache_hit ? _GEN_1821 : dirty_28; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2851 = cache_hit ? _GEN_1822 : dirty_29; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2852 = cache_hit ? _GEN_1823 : dirty_30; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2853 = cache_hit ? _GEN_1824 : dirty_31; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2854 = cache_hit ? _GEN_1825 : dirty_32; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2855 = cache_hit ? _GEN_1826 : dirty_33; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2856 = cache_hit ? _GEN_1827 : dirty_34; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2857 = cache_hit ? _GEN_1828 : dirty_35; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2858 = cache_hit ? _GEN_1829 : dirty_36; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2859 = cache_hit ? _GEN_1830 : dirty_37; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2860 = cache_hit ? _GEN_1831 : dirty_38; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2861 = cache_hit ? _GEN_1832 : dirty_39; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2862 = cache_hit ? _GEN_1833 : dirty_40; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2863 = cache_hit ? _GEN_1834 : dirty_41; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2864 = cache_hit ? _GEN_1835 : dirty_42; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2865 = cache_hit ? _GEN_1836 : dirty_43; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2866 = cache_hit ? _GEN_1837 : dirty_44; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2867 = cache_hit ? _GEN_1838 : dirty_45; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2868 = cache_hit ? _GEN_1839 : dirty_46; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2869 = cache_hit ? _GEN_1840 : dirty_47; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2870 = cache_hit ? _GEN_1841 : dirty_48; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2871 = cache_hit ? _GEN_1842 : dirty_49; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2872 = cache_hit ? _GEN_1843 : dirty_50; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2873 = cache_hit ? _GEN_1844 : dirty_51; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2874 = cache_hit ? _GEN_1845 : dirty_52; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2875 = cache_hit ? _GEN_1846 : dirty_53; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2876 = cache_hit ? _GEN_1847 : dirty_54; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2877 = cache_hit ? _GEN_1848 : dirty_55; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2878 = cache_hit ? _GEN_1849 : dirty_56; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2879 = cache_hit ? _GEN_1850 : dirty_57; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2880 = cache_hit ? _GEN_1851 : dirty_58; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2881 = cache_hit ? _GEN_1852 : dirty_59; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2882 = cache_hit ? _GEN_1853 : dirty_60; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2883 = cache_hit ? _GEN_1854 : dirty_61; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2884 = cache_hit ? _GEN_1855 : dirty_62; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2885 = cache_hit ? _GEN_1856 : dirty_63; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2886 = cache_hit ? _GEN_1857 : dirty_64; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2887 = cache_hit ? _GEN_1858 : dirty_65; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2888 = cache_hit ? _GEN_1859 : dirty_66; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2889 = cache_hit ? _GEN_1860 : dirty_67; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2890 = cache_hit ? _GEN_1861 : dirty_68; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2891 = cache_hit ? _GEN_1862 : dirty_69; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2892 = cache_hit ? _GEN_1863 : dirty_70; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2893 = cache_hit ? _GEN_1864 : dirty_71; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2894 = cache_hit ? _GEN_1865 : dirty_72; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2895 = cache_hit ? _GEN_1866 : dirty_73; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2896 = cache_hit ? _GEN_1867 : dirty_74; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2897 = cache_hit ? _GEN_1868 : dirty_75; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2898 = cache_hit ? _GEN_1869 : dirty_76; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2899 = cache_hit ? _GEN_1870 : dirty_77; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2900 = cache_hit ? _GEN_1871 : dirty_78; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2901 = cache_hit ? _GEN_1872 : dirty_79; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2902 = cache_hit ? _GEN_1873 : dirty_80; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2903 = cache_hit ? _GEN_1874 : dirty_81; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2904 = cache_hit ? _GEN_1875 : dirty_82; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2905 = cache_hit ? _GEN_1876 : dirty_83; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2906 = cache_hit ? _GEN_1877 : dirty_84; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2907 = cache_hit ? _GEN_1878 : dirty_85; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2908 = cache_hit ? _GEN_1879 : dirty_86; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2909 = cache_hit ? _GEN_1880 : dirty_87; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2910 = cache_hit ? _GEN_1881 : dirty_88; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2911 = cache_hit ? _GEN_1882 : dirty_89; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2912 = cache_hit ? _GEN_1883 : dirty_90; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2913 = cache_hit ? _GEN_1884 : dirty_91; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2914 = cache_hit ? _GEN_1885 : dirty_92; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2915 = cache_hit ? _GEN_1886 : dirty_93; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2916 = cache_hit ? _GEN_1887 : dirty_94; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2917 = cache_hit ? _GEN_1888 : dirty_95; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2918 = cache_hit ? _GEN_1889 : dirty_96; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2919 = cache_hit ? _GEN_1890 : dirty_97; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2920 = cache_hit ? _GEN_1891 : dirty_98; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2921 = cache_hit ? _GEN_1892 : dirty_99; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2922 = cache_hit ? _GEN_1893 : dirty_100; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2923 = cache_hit ? _GEN_1894 : dirty_101; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2924 = cache_hit ? _GEN_1895 : dirty_102; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2925 = cache_hit ? _GEN_1896 : dirty_103; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2926 = cache_hit ? _GEN_1897 : dirty_104; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2927 = cache_hit ? _GEN_1898 : dirty_105; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2928 = cache_hit ? _GEN_1899 : dirty_106; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2929 = cache_hit ? _GEN_1900 : dirty_107; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2930 = cache_hit ? _GEN_1901 : dirty_108; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2931 = cache_hit ? _GEN_1902 : dirty_109; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2932 = cache_hit ? _GEN_1903 : dirty_110; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2933 = cache_hit ? _GEN_1904 : dirty_111; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2934 = cache_hit ? _GEN_1905 : dirty_112; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2935 = cache_hit ? _GEN_1906 : dirty_113; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2936 = cache_hit ? _GEN_1907 : dirty_114; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2937 = cache_hit ? _GEN_1908 : dirty_115; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2938 = cache_hit ? _GEN_1909 : dirty_116; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2939 = cache_hit ? _GEN_1910 : dirty_117; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2940 = cache_hit ? _GEN_1911 : dirty_118; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2941 = cache_hit ? _GEN_1912 : dirty_119; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2942 = cache_hit ? _GEN_1913 : dirty_120; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2943 = cache_hit ? _GEN_1914 : dirty_121; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2944 = cache_hit ? _GEN_1915 : dirty_122; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2945 = cache_hit ? _GEN_1916 : dirty_123; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2946 = cache_hit ? _GEN_1917 : dirty_124; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2947 = cache_hit ? _GEN_1918 : dirty_125; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2948 = cache_hit ? _GEN_1919 : dirty_126; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2949 = cache_hit ? _GEN_1920 : dirty_127; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2950 = cache_hit ? _GEN_1921 : dirty_128; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2951 = cache_hit ? _GEN_1922 : dirty_129; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2952 = cache_hit ? _GEN_1923 : dirty_130; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2953 = cache_hit ? _GEN_1924 : dirty_131; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2954 = cache_hit ? _GEN_1925 : dirty_132; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2955 = cache_hit ? _GEN_1926 : dirty_133; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2956 = cache_hit ? _GEN_1927 : dirty_134; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2957 = cache_hit ? _GEN_1928 : dirty_135; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2958 = cache_hit ? _GEN_1929 : dirty_136; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2959 = cache_hit ? _GEN_1930 : dirty_137; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2960 = cache_hit ? _GEN_1931 : dirty_138; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2961 = cache_hit ? _GEN_1932 : dirty_139; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2962 = cache_hit ? _GEN_1933 : dirty_140; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2963 = cache_hit ? _GEN_1934 : dirty_141; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2964 = cache_hit ? _GEN_1935 : dirty_142; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2965 = cache_hit ? _GEN_1936 : dirty_143; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2966 = cache_hit ? _GEN_1937 : dirty_144; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2967 = cache_hit ? _GEN_1938 : dirty_145; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2968 = cache_hit ? _GEN_1939 : dirty_146; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2969 = cache_hit ? _GEN_1940 : dirty_147; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2970 = cache_hit ? _GEN_1941 : dirty_148; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2971 = cache_hit ? _GEN_1942 : dirty_149; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2972 = cache_hit ? _GEN_1943 : dirty_150; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2973 = cache_hit ? _GEN_1944 : dirty_151; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2974 = cache_hit ? _GEN_1945 : dirty_152; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2975 = cache_hit ? _GEN_1946 : dirty_153; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2976 = cache_hit ? _GEN_1947 : dirty_154; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2977 = cache_hit ? _GEN_1948 : dirty_155; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2978 = cache_hit ? _GEN_1949 : dirty_156; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2979 = cache_hit ? _GEN_1950 : dirty_157; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2980 = cache_hit ? _GEN_1951 : dirty_158; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2981 = cache_hit ? _GEN_1952 : dirty_159; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2982 = cache_hit ? _GEN_1953 : dirty_160; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2983 = cache_hit ? _GEN_1954 : dirty_161; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2984 = cache_hit ? _GEN_1955 : dirty_162; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2985 = cache_hit ? _GEN_1956 : dirty_163; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2986 = cache_hit ? _GEN_1957 : dirty_164; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2987 = cache_hit ? _GEN_1958 : dirty_165; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2988 = cache_hit ? _GEN_1959 : dirty_166; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2989 = cache_hit ? _GEN_1960 : dirty_167; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2990 = cache_hit ? _GEN_1961 : dirty_168; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2991 = cache_hit ? _GEN_1962 : dirty_169; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2992 = cache_hit ? _GEN_1963 : dirty_170; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2993 = cache_hit ? _GEN_1964 : dirty_171; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2994 = cache_hit ? _GEN_1965 : dirty_172; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2995 = cache_hit ? _GEN_1966 : dirty_173; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2996 = cache_hit ? _GEN_1967 : dirty_174; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2997 = cache_hit ? _GEN_1968 : dirty_175; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2998 = cache_hit ? _GEN_1969 : dirty_176; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_2999 = cache_hit ? _GEN_1970 : dirty_177; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3000 = cache_hit ? _GEN_1971 : dirty_178; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3001 = cache_hit ? _GEN_1972 : dirty_179; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3002 = cache_hit ? _GEN_1973 : dirty_180; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3003 = cache_hit ? _GEN_1974 : dirty_181; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3004 = cache_hit ? _GEN_1975 : dirty_182; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3005 = cache_hit ? _GEN_1976 : dirty_183; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3006 = cache_hit ? _GEN_1977 : dirty_184; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3007 = cache_hit ? _GEN_1978 : dirty_185; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3008 = cache_hit ? _GEN_1979 : dirty_186; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3009 = cache_hit ? _GEN_1980 : dirty_187; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3010 = cache_hit ? _GEN_1981 : dirty_188; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3011 = cache_hit ? _GEN_1982 : dirty_189; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3012 = cache_hit ? _GEN_1983 : dirty_190; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3013 = cache_hit ? _GEN_1984 : dirty_191; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3014 = cache_hit ? _GEN_1985 : dirty_192; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3015 = cache_hit ? _GEN_1986 : dirty_193; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3016 = cache_hit ? _GEN_1987 : dirty_194; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3017 = cache_hit ? _GEN_1988 : dirty_195; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3018 = cache_hit ? _GEN_1989 : dirty_196; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3019 = cache_hit ? _GEN_1990 : dirty_197; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3020 = cache_hit ? _GEN_1991 : dirty_198; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3021 = cache_hit ? _GEN_1992 : dirty_199; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3022 = cache_hit ? _GEN_1993 : dirty_200; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3023 = cache_hit ? _GEN_1994 : dirty_201; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3024 = cache_hit ? _GEN_1995 : dirty_202; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3025 = cache_hit ? _GEN_1996 : dirty_203; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3026 = cache_hit ? _GEN_1997 : dirty_204; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3027 = cache_hit ? _GEN_1998 : dirty_205; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3028 = cache_hit ? _GEN_1999 : dirty_206; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3029 = cache_hit ? _GEN_2000 : dirty_207; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3030 = cache_hit ? _GEN_2001 : dirty_208; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3031 = cache_hit ? _GEN_2002 : dirty_209; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3032 = cache_hit ? _GEN_2003 : dirty_210; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3033 = cache_hit ? _GEN_2004 : dirty_211; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3034 = cache_hit ? _GEN_2005 : dirty_212; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3035 = cache_hit ? _GEN_2006 : dirty_213; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3036 = cache_hit ? _GEN_2007 : dirty_214; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3037 = cache_hit ? _GEN_2008 : dirty_215; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3038 = cache_hit ? _GEN_2009 : dirty_216; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3039 = cache_hit ? _GEN_2010 : dirty_217; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3040 = cache_hit ? _GEN_2011 : dirty_218; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3041 = cache_hit ? _GEN_2012 : dirty_219; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3042 = cache_hit ? _GEN_2013 : dirty_220; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3043 = cache_hit ? _GEN_2014 : dirty_221; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3044 = cache_hit ? _GEN_2015 : dirty_222; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3045 = cache_hit ? _GEN_2016 : dirty_223; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3046 = cache_hit ? _GEN_2017 : dirty_224; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3047 = cache_hit ? _GEN_2018 : dirty_225; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3048 = cache_hit ? _GEN_2019 : dirty_226; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3049 = cache_hit ? _GEN_2020 : dirty_227; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3050 = cache_hit ? _GEN_2021 : dirty_228; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3051 = cache_hit ? _GEN_2022 : dirty_229; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3052 = cache_hit ? _GEN_2023 : dirty_230; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3053 = cache_hit ? _GEN_2024 : dirty_231; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3054 = cache_hit ? _GEN_2025 : dirty_232; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3055 = cache_hit ? _GEN_2026 : dirty_233; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3056 = cache_hit ? _GEN_2027 : dirty_234; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3057 = cache_hit ? _GEN_2028 : dirty_235; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3058 = cache_hit ? _GEN_2029 : dirty_236; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3059 = cache_hit ? _GEN_2030 : dirty_237; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3060 = cache_hit ? _GEN_2031 : dirty_238; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3061 = cache_hit ? _GEN_2032 : dirty_239; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3062 = cache_hit ? _GEN_2033 : dirty_240; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3063 = cache_hit ? _GEN_2034 : dirty_241; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3064 = cache_hit ? _GEN_2035 : dirty_242; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3065 = cache_hit ? _GEN_2036 : dirty_243; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3066 = cache_hit ? _GEN_2037 : dirty_244; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3067 = cache_hit ? _GEN_2038 : dirty_245; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3068 = cache_hit ? _GEN_2039 : dirty_246; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3069 = cache_hit ? _GEN_2040 : dirty_247; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3070 = cache_hit ? _GEN_2041 : dirty_248; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3071 = cache_hit ? _GEN_2042 : dirty_249; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3072 = cache_hit ? _GEN_2043 : dirty_250; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3073 = cache_hit ? _GEN_2044 : dirty_251; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3074 = cache_hit ? _GEN_2045 : dirty_252; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3075 = cache_hit ? _GEN_2046 : dirty_253; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3076 = cache_hit ? _GEN_2047 : dirty_254; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire  _GEN_3077 = cache_hit ? _GEN_2048 : dirty_255; // @[Dcache.scala 134:29 Dcache.scala 18:24]
  wire [2:0] _GEN_3078 = cache_hit ? 3'h0 : _GEN_2049; // @[Dcache.scala 134:29 Dcache.scala 145:27]
  wire  _T_4 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_4109 = 8'h1 == req_index ? offset_1 : offset_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4110 = 8'h2 == req_index ? offset_2 : _GEN_4109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4111 = 8'h3 == req_index ? offset_3 : _GEN_4110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4112 = 8'h4 == req_index ? offset_4 : _GEN_4111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4113 = 8'h5 == req_index ? offset_5 : _GEN_4112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4114 = 8'h6 == req_index ? offset_6 : _GEN_4113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4115 = 8'h7 == req_index ? offset_7 : _GEN_4114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4116 = 8'h8 == req_index ? offset_8 : _GEN_4115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4117 = 8'h9 == req_index ? offset_9 : _GEN_4116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4118 = 8'ha == req_index ? offset_10 : _GEN_4117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4119 = 8'hb == req_index ? offset_11 : _GEN_4118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4120 = 8'hc == req_index ? offset_12 : _GEN_4119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4121 = 8'hd == req_index ? offset_13 : _GEN_4120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4122 = 8'he == req_index ? offset_14 : _GEN_4121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4123 = 8'hf == req_index ? offset_15 : _GEN_4122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4124 = 8'h10 == req_index ? offset_16 : _GEN_4123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4125 = 8'h11 == req_index ? offset_17 : _GEN_4124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4126 = 8'h12 == req_index ? offset_18 : _GEN_4125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4127 = 8'h13 == req_index ? offset_19 : _GEN_4126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4128 = 8'h14 == req_index ? offset_20 : _GEN_4127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4129 = 8'h15 == req_index ? offset_21 : _GEN_4128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4130 = 8'h16 == req_index ? offset_22 : _GEN_4129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4131 = 8'h17 == req_index ? offset_23 : _GEN_4130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4132 = 8'h18 == req_index ? offset_24 : _GEN_4131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4133 = 8'h19 == req_index ? offset_25 : _GEN_4132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4134 = 8'h1a == req_index ? offset_26 : _GEN_4133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4135 = 8'h1b == req_index ? offset_27 : _GEN_4134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4136 = 8'h1c == req_index ? offset_28 : _GEN_4135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4137 = 8'h1d == req_index ? offset_29 : _GEN_4136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4138 = 8'h1e == req_index ? offset_30 : _GEN_4137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4139 = 8'h1f == req_index ? offset_31 : _GEN_4138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4140 = 8'h20 == req_index ? offset_32 : _GEN_4139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4141 = 8'h21 == req_index ? offset_33 : _GEN_4140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4142 = 8'h22 == req_index ? offset_34 : _GEN_4141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4143 = 8'h23 == req_index ? offset_35 : _GEN_4142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4144 = 8'h24 == req_index ? offset_36 : _GEN_4143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4145 = 8'h25 == req_index ? offset_37 : _GEN_4144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4146 = 8'h26 == req_index ? offset_38 : _GEN_4145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4147 = 8'h27 == req_index ? offset_39 : _GEN_4146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4148 = 8'h28 == req_index ? offset_40 : _GEN_4147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4149 = 8'h29 == req_index ? offset_41 : _GEN_4148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4150 = 8'h2a == req_index ? offset_42 : _GEN_4149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4151 = 8'h2b == req_index ? offset_43 : _GEN_4150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4152 = 8'h2c == req_index ? offset_44 : _GEN_4151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4153 = 8'h2d == req_index ? offset_45 : _GEN_4152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4154 = 8'h2e == req_index ? offset_46 : _GEN_4153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4155 = 8'h2f == req_index ? offset_47 : _GEN_4154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4156 = 8'h30 == req_index ? offset_48 : _GEN_4155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4157 = 8'h31 == req_index ? offset_49 : _GEN_4156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4158 = 8'h32 == req_index ? offset_50 : _GEN_4157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4159 = 8'h33 == req_index ? offset_51 : _GEN_4158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4160 = 8'h34 == req_index ? offset_52 : _GEN_4159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4161 = 8'h35 == req_index ? offset_53 : _GEN_4160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4162 = 8'h36 == req_index ? offset_54 : _GEN_4161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4163 = 8'h37 == req_index ? offset_55 : _GEN_4162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4164 = 8'h38 == req_index ? offset_56 : _GEN_4163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4165 = 8'h39 == req_index ? offset_57 : _GEN_4164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4166 = 8'h3a == req_index ? offset_58 : _GEN_4165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4167 = 8'h3b == req_index ? offset_59 : _GEN_4166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4168 = 8'h3c == req_index ? offset_60 : _GEN_4167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4169 = 8'h3d == req_index ? offset_61 : _GEN_4168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4170 = 8'h3e == req_index ? offset_62 : _GEN_4169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4171 = 8'h3f == req_index ? offset_63 : _GEN_4170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4172 = 8'h40 == req_index ? offset_64 : _GEN_4171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4173 = 8'h41 == req_index ? offset_65 : _GEN_4172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4174 = 8'h42 == req_index ? offset_66 : _GEN_4173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4175 = 8'h43 == req_index ? offset_67 : _GEN_4174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4176 = 8'h44 == req_index ? offset_68 : _GEN_4175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4177 = 8'h45 == req_index ? offset_69 : _GEN_4176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4178 = 8'h46 == req_index ? offset_70 : _GEN_4177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4179 = 8'h47 == req_index ? offset_71 : _GEN_4178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4180 = 8'h48 == req_index ? offset_72 : _GEN_4179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4181 = 8'h49 == req_index ? offset_73 : _GEN_4180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4182 = 8'h4a == req_index ? offset_74 : _GEN_4181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4183 = 8'h4b == req_index ? offset_75 : _GEN_4182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4184 = 8'h4c == req_index ? offset_76 : _GEN_4183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4185 = 8'h4d == req_index ? offset_77 : _GEN_4184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4186 = 8'h4e == req_index ? offset_78 : _GEN_4185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4187 = 8'h4f == req_index ? offset_79 : _GEN_4186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4188 = 8'h50 == req_index ? offset_80 : _GEN_4187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4189 = 8'h51 == req_index ? offset_81 : _GEN_4188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4190 = 8'h52 == req_index ? offset_82 : _GEN_4189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4191 = 8'h53 == req_index ? offset_83 : _GEN_4190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4192 = 8'h54 == req_index ? offset_84 : _GEN_4191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4193 = 8'h55 == req_index ? offset_85 : _GEN_4192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4194 = 8'h56 == req_index ? offset_86 : _GEN_4193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4195 = 8'h57 == req_index ? offset_87 : _GEN_4194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4196 = 8'h58 == req_index ? offset_88 : _GEN_4195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4197 = 8'h59 == req_index ? offset_89 : _GEN_4196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4198 = 8'h5a == req_index ? offset_90 : _GEN_4197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4199 = 8'h5b == req_index ? offset_91 : _GEN_4198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4200 = 8'h5c == req_index ? offset_92 : _GEN_4199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4201 = 8'h5d == req_index ? offset_93 : _GEN_4200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4202 = 8'h5e == req_index ? offset_94 : _GEN_4201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4203 = 8'h5f == req_index ? offset_95 : _GEN_4202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4204 = 8'h60 == req_index ? offset_96 : _GEN_4203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4205 = 8'h61 == req_index ? offset_97 : _GEN_4204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4206 = 8'h62 == req_index ? offset_98 : _GEN_4205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4207 = 8'h63 == req_index ? offset_99 : _GEN_4206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4208 = 8'h64 == req_index ? offset_100 : _GEN_4207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4209 = 8'h65 == req_index ? offset_101 : _GEN_4208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4210 = 8'h66 == req_index ? offset_102 : _GEN_4209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4211 = 8'h67 == req_index ? offset_103 : _GEN_4210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4212 = 8'h68 == req_index ? offset_104 : _GEN_4211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4213 = 8'h69 == req_index ? offset_105 : _GEN_4212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4214 = 8'h6a == req_index ? offset_106 : _GEN_4213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4215 = 8'h6b == req_index ? offset_107 : _GEN_4214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4216 = 8'h6c == req_index ? offset_108 : _GEN_4215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4217 = 8'h6d == req_index ? offset_109 : _GEN_4216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4218 = 8'h6e == req_index ? offset_110 : _GEN_4217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4219 = 8'h6f == req_index ? offset_111 : _GEN_4218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4220 = 8'h70 == req_index ? offset_112 : _GEN_4219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4221 = 8'h71 == req_index ? offset_113 : _GEN_4220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4222 = 8'h72 == req_index ? offset_114 : _GEN_4221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4223 = 8'h73 == req_index ? offset_115 : _GEN_4222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4224 = 8'h74 == req_index ? offset_116 : _GEN_4223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4225 = 8'h75 == req_index ? offset_117 : _GEN_4224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4226 = 8'h76 == req_index ? offset_118 : _GEN_4225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4227 = 8'h77 == req_index ? offset_119 : _GEN_4226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4228 = 8'h78 == req_index ? offset_120 : _GEN_4227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4229 = 8'h79 == req_index ? offset_121 : _GEN_4228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4230 = 8'h7a == req_index ? offset_122 : _GEN_4229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4231 = 8'h7b == req_index ? offset_123 : _GEN_4230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4232 = 8'h7c == req_index ? offset_124 : _GEN_4231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4233 = 8'h7d == req_index ? offset_125 : _GEN_4232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4234 = 8'h7e == req_index ? offset_126 : _GEN_4233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4235 = 8'h7f == req_index ? offset_127 : _GEN_4234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4236 = 8'h80 == req_index ? offset_128 : _GEN_4235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4237 = 8'h81 == req_index ? offset_129 : _GEN_4236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4238 = 8'h82 == req_index ? offset_130 : _GEN_4237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4239 = 8'h83 == req_index ? offset_131 : _GEN_4238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4240 = 8'h84 == req_index ? offset_132 : _GEN_4239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4241 = 8'h85 == req_index ? offset_133 : _GEN_4240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4242 = 8'h86 == req_index ? offset_134 : _GEN_4241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4243 = 8'h87 == req_index ? offset_135 : _GEN_4242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4244 = 8'h88 == req_index ? offset_136 : _GEN_4243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4245 = 8'h89 == req_index ? offset_137 : _GEN_4244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4246 = 8'h8a == req_index ? offset_138 : _GEN_4245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4247 = 8'h8b == req_index ? offset_139 : _GEN_4246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4248 = 8'h8c == req_index ? offset_140 : _GEN_4247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4249 = 8'h8d == req_index ? offset_141 : _GEN_4248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4250 = 8'h8e == req_index ? offset_142 : _GEN_4249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4251 = 8'h8f == req_index ? offset_143 : _GEN_4250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4252 = 8'h90 == req_index ? offset_144 : _GEN_4251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4253 = 8'h91 == req_index ? offset_145 : _GEN_4252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4254 = 8'h92 == req_index ? offset_146 : _GEN_4253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4255 = 8'h93 == req_index ? offset_147 : _GEN_4254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4256 = 8'h94 == req_index ? offset_148 : _GEN_4255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4257 = 8'h95 == req_index ? offset_149 : _GEN_4256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4258 = 8'h96 == req_index ? offset_150 : _GEN_4257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4259 = 8'h97 == req_index ? offset_151 : _GEN_4258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4260 = 8'h98 == req_index ? offset_152 : _GEN_4259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4261 = 8'h99 == req_index ? offset_153 : _GEN_4260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4262 = 8'h9a == req_index ? offset_154 : _GEN_4261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4263 = 8'h9b == req_index ? offset_155 : _GEN_4262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4264 = 8'h9c == req_index ? offset_156 : _GEN_4263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4265 = 8'h9d == req_index ? offset_157 : _GEN_4264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4266 = 8'h9e == req_index ? offset_158 : _GEN_4265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4267 = 8'h9f == req_index ? offset_159 : _GEN_4266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4268 = 8'ha0 == req_index ? offset_160 : _GEN_4267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4269 = 8'ha1 == req_index ? offset_161 : _GEN_4268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4270 = 8'ha2 == req_index ? offset_162 : _GEN_4269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4271 = 8'ha3 == req_index ? offset_163 : _GEN_4270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4272 = 8'ha4 == req_index ? offset_164 : _GEN_4271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4273 = 8'ha5 == req_index ? offset_165 : _GEN_4272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4274 = 8'ha6 == req_index ? offset_166 : _GEN_4273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4275 = 8'ha7 == req_index ? offset_167 : _GEN_4274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4276 = 8'ha8 == req_index ? offset_168 : _GEN_4275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4277 = 8'ha9 == req_index ? offset_169 : _GEN_4276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4278 = 8'haa == req_index ? offset_170 : _GEN_4277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4279 = 8'hab == req_index ? offset_171 : _GEN_4278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4280 = 8'hac == req_index ? offset_172 : _GEN_4279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4281 = 8'had == req_index ? offset_173 : _GEN_4280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4282 = 8'hae == req_index ? offset_174 : _GEN_4281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4283 = 8'haf == req_index ? offset_175 : _GEN_4282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4284 = 8'hb0 == req_index ? offset_176 : _GEN_4283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4285 = 8'hb1 == req_index ? offset_177 : _GEN_4284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4286 = 8'hb2 == req_index ? offset_178 : _GEN_4285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4287 = 8'hb3 == req_index ? offset_179 : _GEN_4286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4288 = 8'hb4 == req_index ? offset_180 : _GEN_4287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4289 = 8'hb5 == req_index ? offset_181 : _GEN_4288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4290 = 8'hb6 == req_index ? offset_182 : _GEN_4289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4291 = 8'hb7 == req_index ? offset_183 : _GEN_4290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4292 = 8'hb8 == req_index ? offset_184 : _GEN_4291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4293 = 8'hb9 == req_index ? offset_185 : _GEN_4292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4294 = 8'hba == req_index ? offset_186 : _GEN_4293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4295 = 8'hbb == req_index ? offset_187 : _GEN_4294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4296 = 8'hbc == req_index ? offset_188 : _GEN_4295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4297 = 8'hbd == req_index ? offset_189 : _GEN_4296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4298 = 8'hbe == req_index ? offset_190 : _GEN_4297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4299 = 8'hbf == req_index ? offset_191 : _GEN_4298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4300 = 8'hc0 == req_index ? offset_192 : _GEN_4299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4301 = 8'hc1 == req_index ? offset_193 : _GEN_4300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4302 = 8'hc2 == req_index ? offset_194 : _GEN_4301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4303 = 8'hc3 == req_index ? offset_195 : _GEN_4302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4304 = 8'hc4 == req_index ? offset_196 : _GEN_4303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4305 = 8'hc5 == req_index ? offset_197 : _GEN_4304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4306 = 8'hc6 == req_index ? offset_198 : _GEN_4305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4307 = 8'hc7 == req_index ? offset_199 : _GEN_4306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4308 = 8'hc8 == req_index ? offset_200 : _GEN_4307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4309 = 8'hc9 == req_index ? offset_201 : _GEN_4308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4310 = 8'hca == req_index ? offset_202 : _GEN_4309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4311 = 8'hcb == req_index ? offset_203 : _GEN_4310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4312 = 8'hcc == req_index ? offset_204 : _GEN_4311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4313 = 8'hcd == req_index ? offset_205 : _GEN_4312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4314 = 8'hce == req_index ? offset_206 : _GEN_4313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4315 = 8'hcf == req_index ? offset_207 : _GEN_4314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4316 = 8'hd0 == req_index ? offset_208 : _GEN_4315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4317 = 8'hd1 == req_index ? offset_209 : _GEN_4316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4318 = 8'hd2 == req_index ? offset_210 : _GEN_4317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4319 = 8'hd3 == req_index ? offset_211 : _GEN_4318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4320 = 8'hd4 == req_index ? offset_212 : _GEN_4319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4321 = 8'hd5 == req_index ? offset_213 : _GEN_4320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4322 = 8'hd6 == req_index ? offset_214 : _GEN_4321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4323 = 8'hd7 == req_index ? offset_215 : _GEN_4322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4324 = 8'hd8 == req_index ? offset_216 : _GEN_4323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4325 = 8'hd9 == req_index ? offset_217 : _GEN_4324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4326 = 8'hda == req_index ? offset_218 : _GEN_4325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4327 = 8'hdb == req_index ? offset_219 : _GEN_4326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4328 = 8'hdc == req_index ? offset_220 : _GEN_4327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4329 = 8'hdd == req_index ? offset_221 : _GEN_4328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4330 = 8'hde == req_index ? offset_222 : _GEN_4329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4331 = 8'hdf == req_index ? offset_223 : _GEN_4330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4332 = 8'he0 == req_index ? offset_224 : _GEN_4331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4333 = 8'he1 == req_index ? offset_225 : _GEN_4332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4334 = 8'he2 == req_index ? offset_226 : _GEN_4333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4335 = 8'he3 == req_index ? offset_227 : _GEN_4334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4336 = 8'he4 == req_index ? offset_228 : _GEN_4335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4337 = 8'he5 == req_index ? offset_229 : _GEN_4336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4338 = 8'he6 == req_index ? offset_230 : _GEN_4337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4339 = 8'he7 == req_index ? offset_231 : _GEN_4338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4340 = 8'he8 == req_index ? offset_232 : _GEN_4339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4341 = 8'he9 == req_index ? offset_233 : _GEN_4340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4342 = 8'hea == req_index ? offset_234 : _GEN_4341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4343 = 8'heb == req_index ? offset_235 : _GEN_4342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4344 = 8'hec == req_index ? offset_236 : _GEN_4343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4345 = 8'hed == req_index ? offset_237 : _GEN_4344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4346 = 8'hee == req_index ? offset_238 : _GEN_4345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4347 = 8'hef == req_index ? offset_239 : _GEN_4346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4348 = 8'hf0 == req_index ? offset_240 : _GEN_4347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4349 = 8'hf1 == req_index ? offset_241 : _GEN_4348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4350 = 8'hf2 == req_index ? offset_242 : _GEN_4349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4351 = 8'hf3 == req_index ? offset_243 : _GEN_4350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4352 = 8'hf4 == req_index ? offset_244 : _GEN_4351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4353 = 8'hf5 == req_index ? offset_245 : _GEN_4352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4354 = 8'hf6 == req_index ? offset_246 : _GEN_4353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4355 = 8'hf7 == req_index ? offset_247 : _GEN_4354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4356 = 8'hf8 == req_index ? offset_248 : _GEN_4355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4357 = 8'hf9 == req_index ? offset_249 : _GEN_4356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4358 = 8'hfa == req_index ? offset_250 : _GEN_4357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4359 = 8'hfb == req_index ? offset_251 : _GEN_4358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4360 = 8'hfc == req_index ? offset_252 : _GEN_4359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4361 = 8'hfd == req_index ? offset_253 : _GEN_4360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4362 = 8'hfe == req_index ? offset_254 : _GEN_4361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4363 = 8'hff == req_index ? offset_255 : _GEN_4362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _data_addr_T = {_GEN_255,req_index,_GEN_4363}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_4364 = io_out_data_ready ? 3'h3 : 3'h2; // @[Dcache.scala 162:31 Dcache.scala 163:25 Dcache.scala 168:19]
  wire  _GEN_4365 = io_out_data_ready ? 1'h0 : 1'h1; // @[Dcache.scala 162:31 Dcache.scala 164:25 Dcache.scala 160:21]
  wire  _T_5 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_6 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_7 = ~cache_fill; // @[Dcache.scala 177:13]
  wire [2:0] _GEN_4366 = ~cache_fill ? 3'h4 : 3'h5; // @[Dcache.scala 177:26 Dcache.scala 178:21 Dcache.scala 187:15]
  wire [31:0] _GEN_4367 = ~cache_fill ? io_dmem_data_addr : 32'h0; // @[Dcache.scala 177:26 Dcache.scala 179:21]
  wire [127:0] _cache_wdata_T_5 = {valid_wdata,io_out_data_read[63:0]}; // @[Cat.scala 30:58]
  wire [127:0] _cache_wdata_T_6 = {io_out_data_read[127:64],valid_wdata}; // @[Cat.scala 30:58]
  wire [127:0] _cache_wdata_T_7 = req_offset[3] ? _cache_wdata_T_5 : _cache_wdata_T_6; // @[Dcache.scala 192:44]
  wire [127:0] _cache_wdata_T_8 = io_dmem_data_req ? _cache_wdata_T_7 : io_out_data_read; // @[Dcache.scala 192:27]
  wire  _GEN_4373 = io_out_data_ready | cache_fill; // @[Dcache.scala 189:29 Dcache.scala 190:21 Dcache.scala 116:28]
  wire  _GEN_4374 = io_out_data_ready | cache_wen; // @[Dcache.scala 189:29 Dcache.scala 191:21 Dcache.scala 117:28]
  wire [127:0] _GEN_4375 = io_out_data_ready ? _cache_wdata_T_8 : cache_wdata; // @[Dcache.scala 189:29 Dcache.scala 192:21 Dcache.scala 118:28]
  wire [127:0] _GEN_4376 = io_out_data_ready ? 128'hffffffffffffffffffffffffffffffff : cache_strb; // @[Dcache.scala 189:29 Dcache.scala 193:21 Dcache.scala 119:28]
  wire  _GEN_4377 = io_out_data_ready ? 1'h0 : _T_7; // @[Dcache.scala 189:29 Dcache.scala 194:21]
  wire  _T_8 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_5402 = _T_8 ? 1'h0 : cache_fill; // @[Conditional.scala 39:67 Dcache.scala 199:25 Dcache.scala 116:28]
  wire  _GEN_5403 = _T_8 | data_ready; // @[Conditional.scala 39:67 Dcache.scala 200:25 Dcache.scala 46:28]
  wire  _GEN_5404 = _T_8 ? 1'h0 : cache_wen; // @[Conditional.scala 39:67 Dcache.scala 201:25 Dcache.scala 117:28]
  wire  _GEN_5405 = _T_8 ? _GEN_769 : valid_0; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5406 = _T_8 ? _GEN_770 : valid_1; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5407 = _T_8 ? _GEN_771 : valid_2; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5408 = _T_8 ? _GEN_772 : valid_3; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5409 = _T_8 ? _GEN_773 : valid_4; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5410 = _T_8 ? _GEN_774 : valid_5; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5411 = _T_8 ? _GEN_775 : valid_6; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5412 = _T_8 ? _GEN_776 : valid_7; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5413 = _T_8 ? _GEN_777 : valid_8; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5414 = _T_8 ? _GEN_778 : valid_9; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5415 = _T_8 ? _GEN_779 : valid_10; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5416 = _T_8 ? _GEN_780 : valid_11; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5417 = _T_8 ? _GEN_781 : valid_12; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5418 = _T_8 ? _GEN_782 : valid_13; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5419 = _T_8 ? _GEN_783 : valid_14; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5420 = _T_8 ? _GEN_784 : valid_15; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5421 = _T_8 ? _GEN_785 : valid_16; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5422 = _T_8 ? _GEN_786 : valid_17; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5423 = _T_8 ? _GEN_787 : valid_18; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5424 = _T_8 ? _GEN_788 : valid_19; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5425 = _T_8 ? _GEN_789 : valid_20; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5426 = _T_8 ? _GEN_790 : valid_21; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5427 = _T_8 ? _GEN_791 : valid_22; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5428 = _T_8 ? _GEN_792 : valid_23; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5429 = _T_8 ? _GEN_793 : valid_24; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5430 = _T_8 ? _GEN_794 : valid_25; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5431 = _T_8 ? _GEN_795 : valid_26; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5432 = _T_8 ? _GEN_796 : valid_27; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5433 = _T_8 ? _GEN_797 : valid_28; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5434 = _T_8 ? _GEN_798 : valid_29; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5435 = _T_8 ? _GEN_799 : valid_30; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5436 = _T_8 ? _GEN_800 : valid_31; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5437 = _T_8 ? _GEN_801 : valid_32; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5438 = _T_8 ? _GEN_802 : valid_33; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5439 = _T_8 ? _GEN_803 : valid_34; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5440 = _T_8 ? _GEN_804 : valid_35; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5441 = _T_8 ? _GEN_805 : valid_36; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5442 = _T_8 ? _GEN_806 : valid_37; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5443 = _T_8 ? _GEN_807 : valid_38; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5444 = _T_8 ? _GEN_808 : valid_39; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5445 = _T_8 ? _GEN_809 : valid_40; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5446 = _T_8 ? _GEN_810 : valid_41; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5447 = _T_8 ? _GEN_811 : valid_42; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5448 = _T_8 ? _GEN_812 : valid_43; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5449 = _T_8 ? _GEN_813 : valid_44; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5450 = _T_8 ? _GEN_814 : valid_45; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5451 = _T_8 ? _GEN_815 : valid_46; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5452 = _T_8 ? _GEN_816 : valid_47; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5453 = _T_8 ? _GEN_817 : valid_48; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5454 = _T_8 ? _GEN_818 : valid_49; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5455 = _T_8 ? _GEN_819 : valid_50; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5456 = _T_8 ? _GEN_820 : valid_51; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5457 = _T_8 ? _GEN_821 : valid_52; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5458 = _T_8 ? _GEN_822 : valid_53; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5459 = _T_8 ? _GEN_823 : valid_54; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5460 = _T_8 ? _GEN_824 : valid_55; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5461 = _T_8 ? _GEN_825 : valid_56; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5462 = _T_8 ? _GEN_826 : valid_57; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5463 = _T_8 ? _GEN_827 : valid_58; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5464 = _T_8 ? _GEN_828 : valid_59; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5465 = _T_8 ? _GEN_829 : valid_60; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5466 = _T_8 ? _GEN_830 : valid_61; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5467 = _T_8 ? _GEN_831 : valid_62; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5468 = _T_8 ? _GEN_832 : valid_63; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5469 = _T_8 ? _GEN_833 : valid_64; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5470 = _T_8 ? _GEN_834 : valid_65; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5471 = _T_8 ? _GEN_835 : valid_66; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5472 = _T_8 ? _GEN_836 : valid_67; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5473 = _T_8 ? _GEN_837 : valid_68; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5474 = _T_8 ? _GEN_838 : valid_69; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5475 = _T_8 ? _GEN_839 : valid_70; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5476 = _T_8 ? _GEN_840 : valid_71; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5477 = _T_8 ? _GEN_841 : valid_72; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5478 = _T_8 ? _GEN_842 : valid_73; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5479 = _T_8 ? _GEN_843 : valid_74; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5480 = _T_8 ? _GEN_844 : valid_75; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5481 = _T_8 ? _GEN_845 : valid_76; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5482 = _T_8 ? _GEN_846 : valid_77; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5483 = _T_8 ? _GEN_847 : valid_78; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5484 = _T_8 ? _GEN_848 : valid_79; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5485 = _T_8 ? _GEN_849 : valid_80; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5486 = _T_8 ? _GEN_850 : valid_81; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5487 = _T_8 ? _GEN_851 : valid_82; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5488 = _T_8 ? _GEN_852 : valid_83; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5489 = _T_8 ? _GEN_853 : valid_84; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5490 = _T_8 ? _GEN_854 : valid_85; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5491 = _T_8 ? _GEN_855 : valid_86; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5492 = _T_8 ? _GEN_856 : valid_87; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5493 = _T_8 ? _GEN_857 : valid_88; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5494 = _T_8 ? _GEN_858 : valid_89; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5495 = _T_8 ? _GEN_859 : valid_90; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5496 = _T_8 ? _GEN_860 : valid_91; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5497 = _T_8 ? _GEN_861 : valid_92; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5498 = _T_8 ? _GEN_862 : valid_93; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5499 = _T_8 ? _GEN_863 : valid_94; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5500 = _T_8 ? _GEN_864 : valid_95; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5501 = _T_8 ? _GEN_865 : valid_96; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5502 = _T_8 ? _GEN_866 : valid_97; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5503 = _T_8 ? _GEN_867 : valid_98; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5504 = _T_8 ? _GEN_868 : valid_99; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5505 = _T_8 ? _GEN_869 : valid_100; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5506 = _T_8 ? _GEN_870 : valid_101; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5507 = _T_8 ? _GEN_871 : valid_102; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5508 = _T_8 ? _GEN_872 : valid_103; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5509 = _T_8 ? _GEN_873 : valid_104; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5510 = _T_8 ? _GEN_874 : valid_105; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5511 = _T_8 ? _GEN_875 : valid_106; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5512 = _T_8 ? _GEN_876 : valid_107; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5513 = _T_8 ? _GEN_877 : valid_108; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5514 = _T_8 ? _GEN_878 : valid_109; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5515 = _T_8 ? _GEN_879 : valid_110; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5516 = _T_8 ? _GEN_880 : valid_111; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5517 = _T_8 ? _GEN_881 : valid_112; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5518 = _T_8 ? _GEN_882 : valid_113; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5519 = _T_8 ? _GEN_883 : valid_114; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5520 = _T_8 ? _GEN_884 : valid_115; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5521 = _T_8 ? _GEN_885 : valid_116; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5522 = _T_8 ? _GEN_886 : valid_117; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5523 = _T_8 ? _GEN_887 : valid_118; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5524 = _T_8 ? _GEN_888 : valid_119; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5525 = _T_8 ? _GEN_889 : valid_120; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5526 = _T_8 ? _GEN_890 : valid_121; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5527 = _T_8 ? _GEN_891 : valid_122; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5528 = _T_8 ? _GEN_892 : valid_123; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5529 = _T_8 ? _GEN_893 : valid_124; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5530 = _T_8 ? _GEN_894 : valid_125; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5531 = _T_8 ? _GEN_895 : valid_126; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5532 = _T_8 ? _GEN_896 : valid_127; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5533 = _T_8 ? _GEN_897 : valid_128; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5534 = _T_8 ? _GEN_898 : valid_129; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5535 = _T_8 ? _GEN_899 : valid_130; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5536 = _T_8 ? _GEN_900 : valid_131; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5537 = _T_8 ? _GEN_901 : valid_132; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5538 = _T_8 ? _GEN_902 : valid_133; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5539 = _T_8 ? _GEN_903 : valid_134; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5540 = _T_8 ? _GEN_904 : valid_135; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5541 = _T_8 ? _GEN_905 : valid_136; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5542 = _T_8 ? _GEN_906 : valid_137; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5543 = _T_8 ? _GEN_907 : valid_138; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5544 = _T_8 ? _GEN_908 : valid_139; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5545 = _T_8 ? _GEN_909 : valid_140; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5546 = _T_8 ? _GEN_910 : valid_141; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5547 = _T_8 ? _GEN_911 : valid_142; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5548 = _T_8 ? _GEN_912 : valid_143; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5549 = _T_8 ? _GEN_913 : valid_144; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5550 = _T_8 ? _GEN_914 : valid_145; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5551 = _T_8 ? _GEN_915 : valid_146; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5552 = _T_8 ? _GEN_916 : valid_147; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5553 = _T_8 ? _GEN_917 : valid_148; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5554 = _T_8 ? _GEN_918 : valid_149; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5555 = _T_8 ? _GEN_919 : valid_150; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5556 = _T_8 ? _GEN_920 : valid_151; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5557 = _T_8 ? _GEN_921 : valid_152; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5558 = _T_8 ? _GEN_922 : valid_153; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5559 = _T_8 ? _GEN_923 : valid_154; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5560 = _T_8 ? _GEN_924 : valid_155; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5561 = _T_8 ? _GEN_925 : valid_156; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5562 = _T_8 ? _GEN_926 : valid_157; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5563 = _T_8 ? _GEN_927 : valid_158; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5564 = _T_8 ? _GEN_928 : valid_159; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5565 = _T_8 ? _GEN_929 : valid_160; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5566 = _T_8 ? _GEN_930 : valid_161; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5567 = _T_8 ? _GEN_931 : valid_162; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5568 = _T_8 ? _GEN_932 : valid_163; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5569 = _T_8 ? _GEN_933 : valid_164; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5570 = _T_8 ? _GEN_934 : valid_165; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5571 = _T_8 ? _GEN_935 : valid_166; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5572 = _T_8 ? _GEN_936 : valid_167; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5573 = _T_8 ? _GEN_937 : valid_168; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5574 = _T_8 ? _GEN_938 : valid_169; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5575 = _T_8 ? _GEN_939 : valid_170; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5576 = _T_8 ? _GEN_940 : valid_171; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5577 = _T_8 ? _GEN_941 : valid_172; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5578 = _T_8 ? _GEN_942 : valid_173; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5579 = _T_8 ? _GEN_943 : valid_174; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5580 = _T_8 ? _GEN_944 : valid_175; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5581 = _T_8 ? _GEN_945 : valid_176; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5582 = _T_8 ? _GEN_946 : valid_177; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5583 = _T_8 ? _GEN_947 : valid_178; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5584 = _T_8 ? _GEN_948 : valid_179; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5585 = _T_8 ? _GEN_949 : valid_180; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5586 = _T_8 ? _GEN_950 : valid_181; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5587 = _T_8 ? _GEN_951 : valid_182; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5588 = _T_8 ? _GEN_952 : valid_183; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5589 = _T_8 ? _GEN_953 : valid_184; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5590 = _T_8 ? _GEN_954 : valid_185; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5591 = _T_8 ? _GEN_955 : valid_186; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5592 = _T_8 ? _GEN_956 : valid_187; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5593 = _T_8 ? _GEN_957 : valid_188; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5594 = _T_8 ? _GEN_958 : valid_189; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5595 = _T_8 ? _GEN_959 : valid_190; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5596 = _T_8 ? _GEN_960 : valid_191; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5597 = _T_8 ? _GEN_961 : valid_192; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5598 = _T_8 ? _GEN_962 : valid_193; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5599 = _T_8 ? _GEN_963 : valid_194; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5600 = _T_8 ? _GEN_964 : valid_195; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5601 = _T_8 ? _GEN_965 : valid_196; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5602 = _T_8 ? _GEN_966 : valid_197; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5603 = _T_8 ? _GEN_967 : valid_198; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5604 = _T_8 ? _GEN_968 : valid_199; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5605 = _T_8 ? _GEN_969 : valid_200; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5606 = _T_8 ? _GEN_970 : valid_201; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5607 = _T_8 ? _GEN_971 : valid_202; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5608 = _T_8 ? _GEN_972 : valid_203; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5609 = _T_8 ? _GEN_973 : valid_204; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5610 = _T_8 ? _GEN_974 : valid_205; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5611 = _T_8 ? _GEN_975 : valid_206; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5612 = _T_8 ? _GEN_976 : valid_207; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5613 = _T_8 ? _GEN_977 : valid_208; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5614 = _T_8 ? _GEN_978 : valid_209; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5615 = _T_8 ? _GEN_979 : valid_210; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5616 = _T_8 ? _GEN_980 : valid_211; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5617 = _T_8 ? _GEN_981 : valid_212; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5618 = _T_8 ? _GEN_982 : valid_213; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5619 = _T_8 ? _GEN_983 : valid_214; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5620 = _T_8 ? _GEN_984 : valid_215; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5621 = _T_8 ? _GEN_985 : valid_216; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5622 = _T_8 ? _GEN_986 : valid_217; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5623 = _T_8 ? _GEN_987 : valid_218; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5624 = _T_8 ? _GEN_988 : valid_219; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5625 = _T_8 ? _GEN_989 : valid_220; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5626 = _T_8 ? _GEN_990 : valid_221; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5627 = _T_8 ? _GEN_991 : valid_222; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5628 = _T_8 ? _GEN_992 : valid_223; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5629 = _T_8 ? _GEN_993 : valid_224; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5630 = _T_8 ? _GEN_994 : valid_225; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5631 = _T_8 ? _GEN_995 : valid_226; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5632 = _T_8 ? _GEN_996 : valid_227; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5633 = _T_8 ? _GEN_997 : valid_228; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5634 = _T_8 ? _GEN_998 : valid_229; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5635 = _T_8 ? _GEN_999 : valid_230; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5636 = _T_8 ? _GEN_1000 : valid_231; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5637 = _T_8 ? _GEN_1001 : valid_232; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5638 = _T_8 ? _GEN_1002 : valid_233; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5639 = _T_8 ? _GEN_1003 : valid_234; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5640 = _T_8 ? _GEN_1004 : valid_235; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5641 = _T_8 ? _GEN_1005 : valid_236; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5642 = _T_8 ? _GEN_1006 : valid_237; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5643 = _T_8 ? _GEN_1007 : valid_238; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5644 = _T_8 ? _GEN_1008 : valid_239; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5645 = _T_8 ? _GEN_1009 : valid_240; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5646 = _T_8 ? _GEN_1010 : valid_241; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5647 = _T_8 ? _GEN_1011 : valid_242; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5648 = _T_8 ? _GEN_1012 : valid_243; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5649 = _T_8 ? _GEN_1013 : valid_244; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5650 = _T_8 ? _GEN_1014 : valid_245; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5651 = _T_8 ? _GEN_1015 : valid_246; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5652 = _T_8 ? _GEN_1016 : valid_247; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5653 = _T_8 ? _GEN_1017 : valid_248; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5654 = _T_8 ? _GEN_1018 : valid_249; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5655 = _T_8 ? _GEN_1019 : valid_250; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5656 = _T_8 ? _GEN_1020 : valid_251; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5657 = _T_8 ? _GEN_1021 : valid_252; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5658 = _T_8 ? _GEN_1022 : valid_253; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5659 = _T_8 ? _GEN_1023 : valid_254; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5660 = _T_8 ? _GEN_1024 : valid_255; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire [19:0] _GEN_5661 = _T_8 ? _GEN_1025 : tag_0; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5662 = _T_8 ? _GEN_1026 : tag_1; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5663 = _T_8 ? _GEN_1027 : tag_2; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5664 = _T_8 ? _GEN_1028 : tag_3; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5665 = _T_8 ? _GEN_1029 : tag_4; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5666 = _T_8 ? _GEN_1030 : tag_5; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5667 = _T_8 ? _GEN_1031 : tag_6; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5668 = _T_8 ? _GEN_1032 : tag_7; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5669 = _T_8 ? _GEN_1033 : tag_8; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5670 = _T_8 ? _GEN_1034 : tag_9; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5671 = _T_8 ? _GEN_1035 : tag_10; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5672 = _T_8 ? _GEN_1036 : tag_11; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5673 = _T_8 ? _GEN_1037 : tag_12; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5674 = _T_8 ? _GEN_1038 : tag_13; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5675 = _T_8 ? _GEN_1039 : tag_14; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5676 = _T_8 ? _GEN_1040 : tag_15; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5677 = _T_8 ? _GEN_1041 : tag_16; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5678 = _T_8 ? _GEN_1042 : tag_17; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5679 = _T_8 ? _GEN_1043 : tag_18; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5680 = _T_8 ? _GEN_1044 : tag_19; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5681 = _T_8 ? _GEN_1045 : tag_20; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5682 = _T_8 ? _GEN_1046 : tag_21; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5683 = _T_8 ? _GEN_1047 : tag_22; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5684 = _T_8 ? _GEN_1048 : tag_23; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5685 = _T_8 ? _GEN_1049 : tag_24; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5686 = _T_8 ? _GEN_1050 : tag_25; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5687 = _T_8 ? _GEN_1051 : tag_26; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5688 = _T_8 ? _GEN_1052 : tag_27; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5689 = _T_8 ? _GEN_1053 : tag_28; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5690 = _T_8 ? _GEN_1054 : tag_29; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5691 = _T_8 ? _GEN_1055 : tag_30; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5692 = _T_8 ? _GEN_1056 : tag_31; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5693 = _T_8 ? _GEN_1057 : tag_32; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5694 = _T_8 ? _GEN_1058 : tag_33; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5695 = _T_8 ? _GEN_1059 : tag_34; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5696 = _T_8 ? _GEN_1060 : tag_35; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5697 = _T_8 ? _GEN_1061 : tag_36; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5698 = _T_8 ? _GEN_1062 : tag_37; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5699 = _T_8 ? _GEN_1063 : tag_38; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5700 = _T_8 ? _GEN_1064 : tag_39; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5701 = _T_8 ? _GEN_1065 : tag_40; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5702 = _T_8 ? _GEN_1066 : tag_41; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5703 = _T_8 ? _GEN_1067 : tag_42; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5704 = _T_8 ? _GEN_1068 : tag_43; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5705 = _T_8 ? _GEN_1069 : tag_44; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5706 = _T_8 ? _GEN_1070 : tag_45; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5707 = _T_8 ? _GEN_1071 : tag_46; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5708 = _T_8 ? _GEN_1072 : tag_47; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5709 = _T_8 ? _GEN_1073 : tag_48; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5710 = _T_8 ? _GEN_1074 : tag_49; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5711 = _T_8 ? _GEN_1075 : tag_50; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5712 = _T_8 ? _GEN_1076 : tag_51; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5713 = _T_8 ? _GEN_1077 : tag_52; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5714 = _T_8 ? _GEN_1078 : tag_53; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5715 = _T_8 ? _GEN_1079 : tag_54; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5716 = _T_8 ? _GEN_1080 : tag_55; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5717 = _T_8 ? _GEN_1081 : tag_56; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5718 = _T_8 ? _GEN_1082 : tag_57; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5719 = _T_8 ? _GEN_1083 : tag_58; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5720 = _T_8 ? _GEN_1084 : tag_59; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5721 = _T_8 ? _GEN_1085 : tag_60; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5722 = _T_8 ? _GEN_1086 : tag_61; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5723 = _T_8 ? _GEN_1087 : tag_62; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5724 = _T_8 ? _GEN_1088 : tag_63; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5725 = _T_8 ? _GEN_1089 : tag_64; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5726 = _T_8 ? _GEN_1090 : tag_65; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5727 = _T_8 ? _GEN_1091 : tag_66; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5728 = _T_8 ? _GEN_1092 : tag_67; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5729 = _T_8 ? _GEN_1093 : tag_68; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5730 = _T_8 ? _GEN_1094 : tag_69; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5731 = _T_8 ? _GEN_1095 : tag_70; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5732 = _T_8 ? _GEN_1096 : tag_71; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5733 = _T_8 ? _GEN_1097 : tag_72; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5734 = _T_8 ? _GEN_1098 : tag_73; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5735 = _T_8 ? _GEN_1099 : tag_74; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5736 = _T_8 ? _GEN_1100 : tag_75; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5737 = _T_8 ? _GEN_1101 : tag_76; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5738 = _T_8 ? _GEN_1102 : tag_77; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5739 = _T_8 ? _GEN_1103 : tag_78; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5740 = _T_8 ? _GEN_1104 : tag_79; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5741 = _T_8 ? _GEN_1105 : tag_80; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5742 = _T_8 ? _GEN_1106 : tag_81; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5743 = _T_8 ? _GEN_1107 : tag_82; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5744 = _T_8 ? _GEN_1108 : tag_83; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5745 = _T_8 ? _GEN_1109 : tag_84; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5746 = _T_8 ? _GEN_1110 : tag_85; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5747 = _T_8 ? _GEN_1111 : tag_86; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5748 = _T_8 ? _GEN_1112 : tag_87; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5749 = _T_8 ? _GEN_1113 : tag_88; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5750 = _T_8 ? _GEN_1114 : tag_89; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5751 = _T_8 ? _GEN_1115 : tag_90; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5752 = _T_8 ? _GEN_1116 : tag_91; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5753 = _T_8 ? _GEN_1117 : tag_92; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5754 = _T_8 ? _GEN_1118 : tag_93; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5755 = _T_8 ? _GEN_1119 : tag_94; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5756 = _T_8 ? _GEN_1120 : tag_95; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5757 = _T_8 ? _GEN_1121 : tag_96; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5758 = _T_8 ? _GEN_1122 : tag_97; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5759 = _T_8 ? _GEN_1123 : tag_98; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5760 = _T_8 ? _GEN_1124 : tag_99; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5761 = _T_8 ? _GEN_1125 : tag_100; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5762 = _T_8 ? _GEN_1126 : tag_101; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5763 = _T_8 ? _GEN_1127 : tag_102; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5764 = _T_8 ? _GEN_1128 : tag_103; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5765 = _T_8 ? _GEN_1129 : tag_104; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5766 = _T_8 ? _GEN_1130 : tag_105; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5767 = _T_8 ? _GEN_1131 : tag_106; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5768 = _T_8 ? _GEN_1132 : tag_107; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5769 = _T_8 ? _GEN_1133 : tag_108; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5770 = _T_8 ? _GEN_1134 : tag_109; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5771 = _T_8 ? _GEN_1135 : tag_110; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5772 = _T_8 ? _GEN_1136 : tag_111; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5773 = _T_8 ? _GEN_1137 : tag_112; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5774 = _T_8 ? _GEN_1138 : tag_113; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5775 = _T_8 ? _GEN_1139 : tag_114; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5776 = _T_8 ? _GEN_1140 : tag_115; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5777 = _T_8 ? _GEN_1141 : tag_116; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5778 = _T_8 ? _GEN_1142 : tag_117; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5779 = _T_8 ? _GEN_1143 : tag_118; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5780 = _T_8 ? _GEN_1144 : tag_119; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5781 = _T_8 ? _GEN_1145 : tag_120; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5782 = _T_8 ? _GEN_1146 : tag_121; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5783 = _T_8 ? _GEN_1147 : tag_122; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5784 = _T_8 ? _GEN_1148 : tag_123; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5785 = _T_8 ? _GEN_1149 : tag_124; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5786 = _T_8 ? _GEN_1150 : tag_125; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5787 = _T_8 ? _GEN_1151 : tag_126; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5788 = _T_8 ? _GEN_1152 : tag_127; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5789 = _T_8 ? _GEN_1153 : tag_128; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5790 = _T_8 ? _GEN_1154 : tag_129; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5791 = _T_8 ? _GEN_1155 : tag_130; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5792 = _T_8 ? _GEN_1156 : tag_131; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5793 = _T_8 ? _GEN_1157 : tag_132; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5794 = _T_8 ? _GEN_1158 : tag_133; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5795 = _T_8 ? _GEN_1159 : tag_134; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5796 = _T_8 ? _GEN_1160 : tag_135; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5797 = _T_8 ? _GEN_1161 : tag_136; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5798 = _T_8 ? _GEN_1162 : tag_137; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5799 = _T_8 ? _GEN_1163 : tag_138; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5800 = _T_8 ? _GEN_1164 : tag_139; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5801 = _T_8 ? _GEN_1165 : tag_140; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5802 = _T_8 ? _GEN_1166 : tag_141; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5803 = _T_8 ? _GEN_1167 : tag_142; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5804 = _T_8 ? _GEN_1168 : tag_143; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5805 = _T_8 ? _GEN_1169 : tag_144; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5806 = _T_8 ? _GEN_1170 : tag_145; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5807 = _T_8 ? _GEN_1171 : tag_146; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5808 = _T_8 ? _GEN_1172 : tag_147; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5809 = _T_8 ? _GEN_1173 : tag_148; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5810 = _T_8 ? _GEN_1174 : tag_149; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5811 = _T_8 ? _GEN_1175 : tag_150; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5812 = _T_8 ? _GEN_1176 : tag_151; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5813 = _T_8 ? _GEN_1177 : tag_152; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5814 = _T_8 ? _GEN_1178 : tag_153; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5815 = _T_8 ? _GEN_1179 : tag_154; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5816 = _T_8 ? _GEN_1180 : tag_155; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5817 = _T_8 ? _GEN_1181 : tag_156; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5818 = _T_8 ? _GEN_1182 : tag_157; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5819 = _T_8 ? _GEN_1183 : tag_158; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5820 = _T_8 ? _GEN_1184 : tag_159; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5821 = _T_8 ? _GEN_1185 : tag_160; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5822 = _T_8 ? _GEN_1186 : tag_161; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5823 = _T_8 ? _GEN_1187 : tag_162; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5824 = _T_8 ? _GEN_1188 : tag_163; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5825 = _T_8 ? _GEN_1189 : tag_164; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5826 = _T_8 ? _GEN_1190 : tag_165; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5827 = _T_8 ? _GEN_1191 : tag_166; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5828 = _T_8 ? _GEN_1192 : tag_167; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5829 = _T_8 ? _GEN_1193 : tag_168; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5830 = _T_8 ? _GEN_1194 : tag_169; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5831 = _T_8 ? _GEN_1195 : tag_170; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5832 = _T_8 ? _GEN_1196 : tag_171; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5833 = _T_8 ? _GEN_1197 : tag_172; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5834 = _T_8 ? _GEN_1198 : tag_173; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5835 = _T_8 ? _GEN_1199 : tag_174; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5836 = _T_8 ? _GEN_1200 : tag_175; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5837 = _T_8 ? _GEN_1201 : tag_176; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5838 = _T_8 ? _GEN_1202 : tag_177; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5839 = _T_8 ? _GEN_1203 : tag_178; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5840 = _T_8 ? _GEN_1204 : tag_179; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5841 = _T_8 ? _GEN_1205 : tag_180; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5842 = _T_8 ? _GEN_1206 : tag_181; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5843 = _T_8 ? _GEN_1207 : tag_182; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5844 = _T_8 ? _GEN_1208 : tag_183; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5845 = _T_8 ? _GEN_1209 : tag_184; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5846 = _T_8 ? _GEN_1210 : tag_185; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5847 = _T_8 ? _GEN_1211 : tag_186; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5848 = _T_8 ? _GEN_1212 : tag_187; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5849 = _T_8 ? _GEN_1213 : tag_188; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5850 = _T_8 ? _GEN_1214 : tag_189; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5851 = _T_8 ? _GEN_1215 : tag_190; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5852 = _T_8 ? _GEN_1216 : tag_191; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5853 = _T_8 ? _GEN_1217 : tag_192; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5854 = _T_8 ? _GEN_1218 : tag_193; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5855 = _T_8 ? _GEN_1219 : tag_194; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5856 = _T_8 ? _GEN_1220 : tag_195; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5857 = _T_8 ? _GEN_1221 : tag_196; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5858 = _T_8 ? _GEN_1222 : tag_197; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5859 = _T_8 ? _GEN_1223 : tag_198; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5860 = _T_8 ? _GEN_1224 : tag_199; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5861 = _T_8 ? _GEN_1225 : tag_200; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5862 = _T_8 ? _GEN_1226 : tag_201; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5863 = _T_8 ? _GEN_1227 : tag_202; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5864 = _T_8 ? _GEN_1228 : tag_203; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5865 = _T_8 ? _GEN_1229 : tag_204; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5866 = _T_8 ? _GEN_1230 : tag_205; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5867 = _T_8 ? _GEN_1231 : tag_206; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5868 = _T_8 ? _GEN_1232 : tag_207; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5869 = _T_8 ? _GEN_1233 : tag_208; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5870 = _T_8 ? _GEN_1234 : tag_209; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5871 = _T_8 ? _GEN_1235 : tag_210; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5872 = _T_8 ? _GEN_1236 : tag_211; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5873 = _T_8 ? _GEN_1237 : tag_212; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5874 = _T_8 ? _GEN_1238 : tag_213; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5875 = _T_8 ? _GEN_1239 : tag_214; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5876 = _T_8 ? _GEN_1240 : tag_215; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5877 = _T_8 ? _GEN_1241 : tag_216; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5878 = _T_8 ? _GEN_1242 : tag_217; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5879 = _T_8 ? _GEN_1243 : tag_218; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5880 = _T_8 ? _GEN_1244 : tag_219; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5881 = _T_8 ? _GEN_1245 : tag_220; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5882 = _T_8 ? _GEN_1246 : tag_221; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5883 = _T_8 ? _GEN_1247 : tag_222; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5884 = _T_8 ? _GEN_1248 : tag_223; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5885 = _T_8 ? _GEN_1249 : tag_224; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5886 = _T_8 ? _GEN_1250 : tag_225; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5887 = _T_8 ? _GEN_1251 : tag_226; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5888 = _T_8 ? _GEN_1252 : tag_227; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5889 = _T_8 ? _GEN_1253 : tag_228; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5890 = _T_8 ? _GEN_1254 : tag_229; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5891 = _T_8 ? _GEN_1255 : tag_230; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5892 = _T_8 ? _GEN_1256 : tag_231; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5893 = _T_8 ? _GEN_1257 : tag_232; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5894 = _T_8 ? _GEN_1258 : tag_233; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5895 = _T_8 ? _GEN_1259 : tag_234; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5896 = _T_8 ? _GEN_1260 : tag_235; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5897 = _T_8 ? _GEN_1261 : tag_236; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5898 = _T_8 ? _GEN_1262 : tag_237; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5899 = _T_8 ? _GEN_1263 : tag_238; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5900 = _T_8 ? _GEN_1264 : tag_239; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5901 = _T_8 ? _GEN_1265 : tag_240; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5902 = _T_8 ? _GEN_1266 : tag_241; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5903 = _T_8 ? _GEN_1267 : tag_242; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5904 = _T_8 ? _GEN_1268 : tag_243; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5905 = _T_8 ? _GEN_1269 : tag_244; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5906 = _T_8 ? _GEN_1270 : tag_245; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5907 = _T_8 ? _GEN_1271 : tag_246; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5908 = _T_8 ? _GEN_1272 : tag_247; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5909 = _T_8 ? _GEN_1273 : tag_248; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5910 = _T_8 ? _GEN_1274 : tag_249; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5911 = _T_8 ? _GEN_1275 : tag_250; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5912 = _T_8 ? _GEN_1276 : tag_251; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5913 = _T_8 ? _GEN_1277 : tag_252; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5914 = _T_8 ? _GEN_1278 : tag_253; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5915 = _T_8 ? _GEN_1279 : tag_254; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5916 = _T_8 ? _GEN_1280 : tag_255; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire  _GEN_5917 = _T_8 ? _GEN_1537 : dirty_0; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5918 = _T_8 ? _GEN_1538 : dirty_1; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5919 = _T_8 ? _GEN_1539 : dirty_2; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5920 = _T_8 ? _GEN_1540 : dirty_3; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5921 = _T_8 ? _GEN_1541 : dirty_4; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5922 = _T_8 ? _GEN_1542 : dirty_5; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5923 = _T_8 ? _GEN_1543 : dirty_6; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5924 = _T_8 ? _GEN_1544 : dirty_7; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5925 = _T_8 ? _GEN_1545 : dirty_8; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5926 = _T_8 ? _GEN_1546 : dirty_9; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5927 = _T_8 ? _GEN_1547 : dirty_10; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5928 = _T_8 ? _GEN_1548 : dirty_11; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5929 = _T_8 ? _GEN_1549 : dirty_12; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5930 = _T_8 ? _GEN_1550 : dirty_13; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5931 = _T_8 ? _GEN_1551 : dirty_14; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5932 = _T_8 ? _GEN_1552 : dirty_15; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5933 = _T_8 ? _GEN_1553 : dirty_16; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5934 = _T_8 ? _GEN_1554 : dirty_17; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5935 = _T_8 ? _GEN_1555 : dirty_18; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5936 = _T_8 ? _GEN_1556 : dirty_19; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5937 = _T_8 ? _GEN_1557 : dirty_20; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5938 = _T_8 ? _GEN_1558 : dirty_21; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5939 = _T_8 ? _GEN_1559 : dirty_22; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5940 = _T_8 ? _GEN_1560 : dirty_23; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5941 = _T_8 ? _GEN_1561 : dirty_24; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5942 = _T_8 ? _GEN_1562 : dirty_25; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5943 = _T_8 ? _GEN_1563 : dirty_26; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5944 = _T_8 ? _GEN_1564 : dirty_27; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5945 = _T_8 ? _GEN_1565 : dirty_28; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5946 = _T_8 ? _GEN_1566 : dirty_29; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5947 = _T_8 ? _GEN_1567 : dirty_30; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5948 = _T_8 ? _GEN_1568 : dirty_31; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5949 = _T_8 ? _GEN_1569 : dirty_32; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5950 = _T_8 ? _GEN_1570 : dirty_33; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5951 = _T_8 ? _GEN_1571 : dirty_34; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5952 = _T_8 ? _GEN_1572 : dirty_35; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5953 = _T_8 ? _GEN_1573 : dirty_36; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5954 = _T_8 ? _GEN_1574 : dirty_37; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5955 = _T_8 ? _GEN_1575 : dirty_38; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5956 = _T_8 ? _GEN_1576 : dirty_39; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5957 = _T_8 ? _GEN_1577 : dirty_40; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5958 = _T_8 ? _GEN_1578 : dirty_41; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5959 = _T_8 ? _GEN_1579 : dirty_42; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5960 = _T_8 ? _GEN_1580 : dirty_43; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5961 = _T_8 ? _GEN_1581 : dirty_44; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5962 = _T_8 ? _GEN_1582 : dirty_45; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5963 = _T_8 ? _GEN_1583 : dirty_46; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5964 = _T_8 ? _GEN_1584 : dirty_47; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5965 = _T_8 ? _GEN_1585 : dirty_48; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5966 = _T_8 ? _GEN_1586 : dirty_49; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5967 = _T_8 ? _GEN_1587 : dirty_50; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5968 = _T_8 ? _GEN_1588 : dirty_51; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5969 = _T_8 ? _GEN_1589 : dirty_52; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5970 = _T_8 ? _GEN_1590 : dirty_53; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5971 = _T_8 ? _GEN_1591 : dirty_54; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5972 = _T_8 ? _GEN_1592 : dirty_55; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5973 = _T_8 ? _GEN_1593 : dirty_56; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5974 = _T_8 ? _GEN_1594 : dirty_57; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5975 = _T_8 ? _GEN_1595 : dirty_58; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5976 = _T_8 ? _GEN_1596 : dirty_59; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5977 = _T_8 ? _GEN_1597 : dirty_60; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5978 = _T_8 ? _GEN_1598 : dirty_61; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5979 = _T_8 ? _GEN_1599 : dirty_62; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5980 = _T_8 ? _GEN_1600 : dirty_63; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5981 = _T_8 ? _GEN_1601 : dirty_64; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5982 = _T_8 ? _GEN_1602 : dirty_65; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5983 = _T_8 ? _GEN_1603 : dirty_66; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5984 = _T_8 ? _GEN_1604 : dirty_67; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5985 = _T_8 ? _GEN_1605 : dirty_68; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5986 = _T_8 ? _GEN_1606 : dirty_69; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5987 = _T_8 ? _GEN_1607 : dirty_70; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5988 = _T_8 ? _GEN_1608 : dirty_71; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5989 = _T_8 ? _GEN_1609 : dirty_72; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5990 = _T_8 ? _GEN_1610 : dirty_73; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5991 = _T_8 ? _GEN_1611 : dirty_74; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5992 = _T_8 ? _GEN_1612 : dirty_75; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5993 = _T_8 ? _GEN_1613 : dirty_76; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5994 = _T_8 ? _GEN_1614 : dirty_77; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5995 = _T_8 ? _GEN_1615 : dirty_78; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5996 = _T_8 ? _GEN_1616 : dirty_79; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5997 = _T_8 ? _GEN_1617 : dirty_80; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5998 = _T_8 ? _GEN_1618 : dirty_81; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5999 = _T_8 ? _GEN_1619 : dirty_82; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6000 = _T_8 ? _GEN_1620 : dirty_83; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6001 = _T_8 ? _GEN_1621 : dirty_84; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6002 = _T_8 ? _GEN_1622 : dirty_85; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6003 = _T_8 ? _GEN_1623 : dirty_86; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6004 = _T_8 ? _GEN_1624 : dirty_87; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6005 = _T_8 ? _GEN_1625 : dirty_88; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6006 = _T_8 ? _GEN_1626 : dirty_89; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6007 = _T_8 ? _GEN_1627 : dirty_90; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6008 = _T_8 ? _GEN_1628 : dirty_91; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6009 = _T_8 ? _GEN_1629 : dirty_92; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6010 = _T_8 ? _GEN_1630 : dirty_93; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6011 = _T_8 ? _GEN_1631 : dirty_94; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6012 = _T_8 ? _GEN_1632 : dirty_95; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6013 = _T_8 ? _GEN_1633 : dirty_96; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6014 = _T_8 ? _GEN_1634 : dirty_97; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6015 = _T_8 ? _GEN_1635 : dirty_98; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6016 = _T_8 ? _GEN_1636 : dirty_99; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6017 = _T_8 ? _GEN_1637 : dirty_100; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6018 = _T_8 ? _GEN_1638 : dirty_101; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6019 = _T_8 ? _GEN_1639 : dirty_102; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6020 = _T_8 ? _GEN_1640 : dirty_103; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6021 = _T_8 ? _GEN_1641 : dirty_104; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6022 = _T_8 ? _GEN_1642 : dirty_105; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6023 = _T_8 ? _GEN_1643 : dirty_106; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6024 = _T_8 ? _GEN_1644 : dirty_107; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6025 = _T_8 ? _GEN_1645 : dirty_108; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6026 = _T_8 ? _GEN_1646 : dirty_109; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6027 = _T_8 ? _GEN_1647 : dirty_110; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6028 = _T_8 ? _GEN_1648 : dirty_111; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6029 = _T_8 ? _GEN_1649 : dirty_112; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6030 = _T_8 ? _GEN_1650 : dirty_113; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6031 = _T_8 ? _GEN_1651 : dirty_114; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6032 = _T_8 ? _GEN_1652 : dirty_115; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6033 = _T_8 ? _GEN_1653 : dirty_116; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6034 = _T_8 ? _GEN_1654 : dirty_117; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6035 = _T_8 ? _GEN_1655 : dirty_118; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6036 = _T_8 ? _GEN_1656 : dirty_119; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6037 = _T_8 ? _GEN_1657 : dirty_120; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6038 = _T_8 ? _GEN_1658 : dirty_121; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6039 = _T_8 ? _GEN_1659 : dirty_122; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6040 = _T_8 ? _GEN_1660 : dirty_123; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6041 = _T_8 ? _GEN_1661 : dirty_124; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6042 = _T_8 ? _GEN_1662 : dirty_125; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6043 = _T_8 ? _GEN_1663 : dirty_126; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6044 = _T_8 ? _GEN_1664 : dirty_127; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6045 = _T_8 ? _GEN_1665 : dirty_128; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6046 = _T_8 ? _GEN_1666 : dirty_129; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6047 = _T_8 ? _GEN_1667 : dirty_130; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6048 = _T_8 ? _GEN_1668 : dirty_131; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6049 = _T_8 ? _GEN_1669 : dirty_132; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6050 = _T_8 ? _GEN_1670 : dirty_133; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6051 = _T_8 ? _GEN_1671 : dirty_134; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6052 = _T_8 ? _GEN_1672 : dirty_135; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6053 = _T_8 ? _GEN_1673 : dirty_136; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6054 = _T_8 ? _GEN_1674 : dirty_137; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6055 = _T_8 ? _GEN_1675 : dirty_138; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6056 = _T_8 ? _GEN_1676 : dirty_139; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6057 = _T_8 ? _GEN_1677 : dirty_140; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6058 = _T_8 ? _GEN_1678 : dirty_141; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6059 = _T_8 ? _GEN_1679 : dirty_142; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6060 = _T_8 ? _GEN_1680 : dirty_143; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6061 = _T_8 ? _GEN_1681 : dirty_144; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6062 = _T_8 ? _GEN_1682 : dirty_145; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6063 = _T_8 ? _GEN_1683 : dirty_146; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6064 = _T_8 ? _GEN_1684 : dirty_147; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6065 = _T_8 ? _GEN_1685 : dirty_148; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6066 = _T_8 ? _GEN_1686 : dirty_149; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6067 = _T_8 ? _GEN_1687 : dirty_150; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6068 = _T_8 ? _GEN_1688 : dirty_151; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6069 = _T_8 ? _GEN_1689 : dirty_152; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6070 = _T_8 ? _GEN_1690 : dirty_153; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6071 = _T_8 ? _GEN_1691 : dirty_154; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6072 = _T_8 ? _GEN_1692 : dirty_155; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6073 = _T_8 ? _GEN_1693 : dirty_156; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6074 = _T_8 ? _GEN_1694 : dirty_157; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6075 = _T_8 ? _GEN_1695 : dirty_158; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6076 = _T_8 ? _GEN_1696 : dirty_159; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6077 = _T_8 ? _GEN_1697 : dirty_160; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6078 = _T_8 ? _GEN_1698 : dirty_161; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6079 = _T_8 ? _GEN_1699 : dirty_162; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6080 = _T_8 ? _GEN_1700 : dirty_163; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6081 = _T_8 ? _GEN_1701 : dirty_164; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6082 = _T_8 ? _GEN_1702 : dirty_165; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6083 = _T_8 ? _GEN_1703 : dirty_166; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6084 = _T_8 ? _GEN_1704 : dirty_167; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6085 = _T_8 ? _GEN_1705 : dirty_168; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6086 = _T_8 ? _GEN_1706 : dirty_169; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6087 = _T_8 ? _GEN_1707 : dirty_170; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6088 = _T_8 ? _GEN_1708 : dirty_171; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6089 = _T_8 ? _GEN_1709 : dirty_172; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6090 = _T_8 ? _GEN_1710 : dirty_173; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6091 = _T_8 ? _GEN_1711 : dirty_174; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6092 = _T_8 ? _GEN_1712 : dirty_175; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6093 = _T_8 ? _GEN_1713 : dirty_176; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6094 = _T_8 ? _GEN_1714 : dirty_177; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6095 = _T_8 ? _GEN_1715 : dirty_178; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6096 = _T_8 ? _GEN_1716 : dirty_179; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6097 = _T_8 ? _GEN_1717 : dirty_180; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6098 = _T_8 ? _GEN_1718 : dirty_181; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6099 = _T_8 ? _GEN_1719 : dirty_182; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6100 = _T_8 ? _GEN_1720 : dirty_183; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6101 = _T_8 ? _GEN_1721 : dirty_184; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6102 = _T_8 ? _GEN_1722 : dirty_185; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6103 = _T_8 ? _GEN_1723 : dirty_186; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6104 = _T_8 ? _GEN_1724 : dirty_187; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6105 = _T_8 ? _GEN_1725 : dirty_188; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6106 = _T_8 ? _GEN_1726 : dirty_189; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6107 = _T_8 ? _GEN_1727 : dirty_190; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6108 = _T_8 ? _GEN_1728 : dirty_191; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6109 = _T_8 ? _GEN_1729 : dirty_192; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6110 = _T_8 ? _GEN_1730 : dirty_193; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6111 = _T_8 ? _GEN_1731 : dirty_194; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6112 = _T_8 ? _GEN_1732 : dirty_195; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6113 = _T_8 ? _GEN_1733 : dirty_196; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6114 = _T_8 ? _GEN_1734 : dirty_197; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6115 = _T_8 ? _GEN_1735 : dirty_198; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6116 = _T_8 ? _GEN_1736 : dirty_199; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6117 = _T_8 ? _GEN_1737 : dirty_200; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6118 = _T_8 ? _GEN_1738 : dirty_201; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6119 = _T_8 ? _GEN_1739 : dirty_202; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6120 = _T_8 ? _GEN_1740 : dirty_203; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6121 = _T_8 ? _GEN_1741 : dirty_204; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6122 = _T_8 ? _GEN_1742 : dirty_205; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6123 = _T_8 ? _GEN_1743 : dirty_206; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6124 = _T_8 ? _GEN_1744 : dirty_207; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6125 = _T_8 ? _GEN_1745 : dirty_208; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6126 = _T_8 ? _GEN_1746 : dirty_209; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6127 = _T_8 ? _GEN_1747 : dirty_210; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6128 = _T_8 ? _GEN_1748 : dirty_211; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6129 = _T_8 ? _GEN_1749 : dirty_212; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6130 = _T_8 ? _GEN_1750 : dirty_213; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6131 = _T_8 ? _GEN_1751 : dirty_214; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6132 = _T_8 ? _GEN_1752 : dirty_215; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6133 = _T_8 ? _GEN_1753 : dirty_216; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6134 = _T_8 ? _GEN_1754 : dirty_217; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6135 = _T_8 ? _GEN_1755 : dirty_218; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6136 = _T_8 ? _GEN_1756 : dirty_219; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6137 = _T_8 ? _GEN_1757 : dirty_220; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6138 = _T_8 ? _GEN_1758 : dirty_221; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6139 = _T_8 ? _GEN_1759 : dirty_222; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6140 = _T_8 ? _GEN_1760 : dirty_223; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6141 = _T_8 ? _GEN_1761 : dirty_224; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6142 = _T_8 ? _GEN_1762 : dirty_225; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6143 = _T_8 ? _GEN_1763 : dirty_226; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6144 = _T_8 ? _GEN_1764 : dirty_227; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6145 = _T_8 ? _GEN_1765 : dirty_228; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6146 = _T_8 ? _GEN_1766 : dirty_229; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6147 = _T_8 ? _GEN_1767 : dirty_230; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6148 = _T_8 ? _GEN_1768 : dirty_231; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6149 = _T_8 ? _GEN_1769 : dirty_232; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6150 = _T_8 ? _GEN_1770 : dirty_233; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6151 = _T_8 ? _GEN_1771 : dirty_234; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6152 = _T_8 ? _GEN_1772 : dirty_235; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6153 = _T_8 ? _GEN_1773 : dirty_236; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6154 = _T_8 ? _GEN_1774 : dirty_237; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6155 = _T_8 ? _GEN_1775 : dirty_238; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6156 = _T_8 ? _GEN_1776 : dirty_239; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6157 = _T_8 ? _GEN_1777 : dirty_240; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6158 = _T_8 ? _GEN_1778 : dirty_241; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6159 = _T_8 ? _GEN_1779 : dirty_242; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6160 = _T_8 ? _GEN_1780 : dirty_243; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6161 = _T_8 ? _GEN_1781 : dirty_244; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6162 = _T_8 ? _GEN_1782 : dirty_245; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6163 = _T_8 ? _GEN_1783 : dirty_246; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6164 = _T_8 ? _GEN_1784 : dirty_247; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6165 = _T_8 ? _GEN_1785 : dirty_248; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6166 = _T_8 ? _GEN_1786 : dirty_249; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6167 = _T_8 ? _GEN_1787 : dirty_250; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6168 = _T_8 ? _GEN_1788 : dirty_251; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6169 = _T_8 ? _GEN_1789 : dirty_252; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6170 = _T_8 ? _GEN_1790 : dirty_253; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6171 = _T_8 ? _GEN_1791 : dirty_254; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6172 = _T_8 ? _GEN_1792 : dirty_255; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire [3:0] _GEN_6173 = _T_8 ? _GEN_1281 : offset_0; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6174 = _T_8 ? _GEN_1282 : offset_1; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6175 = _T_8 ? _GEN_1283 : offset_2; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6176 = _T_8 ? _GEN_1284 : offset_3; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6177 = _T_8 ? _GEN_1285 : offset_4; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6178 = _T_8 ? _GEN_1286 : offset_5; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6179 = _T_8 ? _GEN_1287 : offset_6; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6180 = _T_8 ? _GEN_1288 : offset_7; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6181 = _T_8 ? _GEN_1289 : offset_8; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6182 = _T_8 ? _GEN_1290 : offset_9; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6183 = _T_8 ? _GEN_1291 : offset_10; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6184 = _T_8 ? _GEN_1292 : offset_11; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6185 = _T_8 ? _GEN_1293 : offset_12; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6186 = _T_8 ? _GEN_1294 : offset_13; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6187 = _T_8 ? _GEN_1295 : offset_14; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6188 = _T_8 ? _GEN_1296 : offset_15; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6189 = _T_8 ? _GEN_1297 : offset_16; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6190 = _T_8 ? _GEN_1298 : offset_17; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6191 = _T_8 ? _GEN_1299 : offset_18; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6192 = _T_8 ? _GEN_1300 : offset_19; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6193 = _T_8 ? _GEN_1301 : offset_20; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6194 = _T_8 ? _GEN_1302 : offset_21; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6195 = _T_8 ? _GEN_1303 : offset_22; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6196 = _T_8 ? _GEN_1304 : offset_23; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6197 = _T_8 ? _GEN_1305 : offset_24; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6198 = _T_8 ? _GEN_1306 : offset_25; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6199 = _T_8 ? _GEN_1307 : offset_26; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6200 = _T_8 ? _GEN_1308 : offset_27; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6201 = _T_8 ? _GEN_1309 : offset_28; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6202 = _T_8 ? _GEN_1310 : offset_29; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6203 = _T_8 ? _GEN_1311 : offset_30; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6204 = _T_8 ? _GEN_1312 : offset_31; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6205 = _T_8 ? _GEN_1313 : offset_32; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6206 = _T_8 ? _GEN_1314 : offset_33; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6207 = _T_8 ? _GEN_1315 : offset_34; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6208 = _T_8 ? _GEN_1316 : offset_35; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6209 = _T_8 ? _GEN_1317 : offset_36; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6210 = _T_8 ? _GEN_1318 : offset_37; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6211 = _T_8 ? _GEN_1319 : offset_38; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6212 = _T_8 ? _GEN_1320 : offset_39; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6213 = _T_8 ? _GEN_1321 : offset_40; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6214 = _T_8 ? _GEN_1322 : offset_41; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6215 = _T_8 ? _GEN_1323 : offset_42; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6216 = _T_8 ? _GEN_1324 : offset_43; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6217 = _T_8 ? _GEN_1325 : offset_44; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6218 = _T_8 ? _GEN_1326 : offset_45; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6219 = _T_8 ? _GEN_1327 : offset_46; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6220 = _T_8 ? _GEN_1328 : offset_47; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6221 = _T_8 ? _GEN_1329 : offset_48; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6222 = _T_8 ? _GEN_1330 : offset_49; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6223 = _T_8 ? _GEN_1331 : offset_50; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6224 = _T_8 ? _GEN_1332 : offset_51; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6225 = _T_8 ? _GEN_1333 : offset_52; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6226 = _T_8 ? _GEN_1334 : offset_53; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6227 = _T_8 ? _GEN_1335 : offset_54; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6228 = _T_8 ? _GEN_1336 : offset_55; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6229 = _T_8 ? _GEN_1337 : offset_56; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6230 = _T_8 ? _GEN_1338 : offset_57; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6231 = _T_8 ? _GEN_1339 : offset_58; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6232 = _T_8 ? _GEN_1340 : offset_59; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6233 = _T_8 ? _GEN_1341 : offset_60; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6234 = _T_8 ? _GEN_1342 : offset_61; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6235 = _T_8 ? _GEN_1343 : offset_62; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6236 = _T_8 ? _GEN_1344 : offset_63; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6237 = _T_8 ? _GEN_1345 : offset_64; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6238 = _T_8 ? _GEN_1346 : offset_65; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6239 = _T_8 ? _GEN_1347 : offset_66; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6240 = _T_8 ? _GEN_1348 : offset_67; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6241 = _T_8 ? _GEN_1349 : offset_68; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6242 = _T_8 ? _GEN_1350 : offset_69; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6243 = _T_8 ? _GEN_1351 : offset_70; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6244 = _T_8 ? _GEN_1352 : offset_71; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6245 = _T_8 ? _GEN_1353 : offset_72; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6246 = _T_8 ? _GEN_1354 : offset_73; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6247 = _T_8 ? _GEN_1355 : offset_74; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6248 = _T_8 ? _GEN_1356 : offset_75; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6249 = _T_8 ? _GEN_1357 : offset_76; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6250 = _T_8 ? _GEN_1358 : offset_77; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6251 = _T_8 ? _GEN_1359 : offset_78; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6252 = _T_8 ? _GEN_1360 : offset_79; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6253 = _T_8 ? _GEN_1361 : offset_80; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6254 = _T_8 ? _GEN_1362 : offset_81; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6255 = _T_8 ? _GEN_1363 : offset_82; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6256 = _T_8 ? _GEN_1364 : offset_83; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6257 = _T_8 ? _GEN_1365 : offset_84; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6258 = _T_8 ? _GEN_1366 : offset_85; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6259 = _T_8 ? _GEN_1367 : offset_86; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6260 = _T_8 ? _GEN_1368 : offset_87; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6261 = _T_8 ? _GEN_1369 : offset_88; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6262 = _T_8 ? _GEN_1370 : offset_89; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6263 = _T_8 ? _GEN_1371 : offset_90; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6264 = _T_8 ? _GEN_1372 : offset_91; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6265 = _T_8 ? _GEN_1373 : offset_92; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6266 = _T_8 ? _GEN_1374 : offset_93; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6267 = _T_8 ? _GEN_1375 : offset_94; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6268 = _T_8 ? _GEN_1376 : offset_95; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6269 = _T_8 ? _GEN_1377 : offset_96; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6270 = _T_8 ? _GEN_1378 : offset_97; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6271 = _T_8 ? _GEN_1379 : offset_98; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6272 = _T_8 ? _GEN_1380 : offset_99; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6273 = _T_8 ? _GEN_1381 : offset_100; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6274 = _T_8 ? _GEN_1382 : offset_101; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6275 = _T_8 ? _GEN_1383 : offset_102; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6276 = _T_8 ? _GEN_1384 : offset_103; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6277 = _T_8 ? _GEN_1385 : offset_104; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6278 = _T_8 ? _GEN_1386 : offset_105; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6279 = _T_8 ? _GEN_1387 : offset_106; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6280 = _T_8 ? _GEN_1388 : offset_107; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6281 = _T_8 ? _GEN_1389 : offset_108; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6282 = _T_8 ? _GEN_1390 : offset_109; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6283 = _T_8 ? _GEN_1391 : offset_110; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6284 = _T_8 ? _GEN_1392 : offset_111; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6285 = _T_8 ? _GEN_1393 : offset_112; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6286 = _T_8 ? _GEN_1394 : offset_113; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6287 = _T_8 ? _GEN_1395 : offset_114; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6288 = _T_8 ? _GEN_1396 : offset_115; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6289 = _T_8 ? _GEN_1397 : offset_116; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6290 = _T_8 ? _GEN_1398 : offset_117; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6291 = _T_8 ? _GEN_1399 : offset_118; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6292 = _T_8 ? _GEN_1400 : offset_119; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6293 = _T_8 ? _GEN_1401 : offset_120; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6294 = _T_8 ? _GEN_1402 : offset_121; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6295 = _T_8 ? _GEN_1403 : offset_122; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6296 = _T_8 ? _GEN_1404 : offset_123; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6297 = _T_8 ? _GEN_1405 : offset_124; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6298 = _T_8 ? _GEN_1406 : offset_125; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6299 = _T_8 ? _GEN_1407 : offset_126; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6300 = _T_8 ? _GEN_1408 : offset_127; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6301 = _T_8 ? _GEN_1409 : offset_128; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6302 = _T_8 ? _GEN_1410 : offset_129; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6303 = _T_8 ? _GEN_1411 : offset_130; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6304 = _T_8 ? _GEN_1412 : offset_131; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6305 = _T_8 ? _GEN_1413 : offset_132; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6306 = _T_8 ? _GEN_1414 : offset_133; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6307 = _T_8 ? _GEN_1415 : offset_134; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6308 = _T_8 ? _GEN_1416 : offset_135; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6309 = _T_8 ? _GEN_1417 : offset_136; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6310 = _T_8 ? _GEN_1418 : offset_137; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6311 = _T_8 ? _GEN_1419 : offset_138; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6312 = _T_8 ? _GEN_1420 : offset_139; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6313 = _T_8 ? _GEN_1421 : offset_140; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6314 = _T_8 ? _GEN_1422 : offset_141; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6315 = _T_8 ? _GEN_1423 : offset_142; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6316 = _T_8 ? _GEN_1424 : offset_143; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6317 = _T_8 ? _GEN_1425 : offset_144; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6318 = _T_8 ? _GEN_1426 : offset_145; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6319 = _T_8 ? _GEN_1427 : offset_146; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6320 = _T_8 ? _GEN_1428 : offset_147; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6321 = _T_8 ? _GEN_1429 : offset_148; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6322 = _T_8 ? _GEN_1430 : offset_149; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6323 = _T_8 ? _GEN_1431 : offset_150; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6324 = _T_8 ? _GEN_1432 : offset_151; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6325 = _T_8 ? _GEN_1433 : offset_152; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6326 = _T_8 ? _GEN_1434 : offset_153; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6327 = _T_8 ? _GEN_1435 : offset_154; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6328 = _T_8 ? _GEN_1436 : offset_155; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6329 = _T_8 ? _GEN_1437 : offset_156; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6330 = _T_8 ? _GEN_1438 : offset_157; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6331 = _T_8 ? _GEN_1439 : offset_158; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6332 = _T_8 ? _GEN_1440 : offset_159; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6333 = _T_8 ? _GEN_1441 : offset_160; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6334 = _T_8 ? _GEN_1442 : offset_161; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6335 = _T_8 ? _GEN_1443 : offset_162; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6336 = _T_8 ? _GEN_1444 : offset_163; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6337 = _T_8 ? _GEN_1445 : offset_164; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6338 = _T_8 ? _GEN_1446 : offset_165; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6339 = _T_8 ? _GEN_1447 : offset_166; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6340 = _T_8 ? _GEN_1448 : offset_167; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6341 = _T_8 ? _GEN_1449 : offset_168; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6342 = _T_8 ? _GEN_1450 : offset_169; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6343 = _T_8 ? _GEN_1451 : offset_170; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6344 = _T_8 ? _GEN_1452 : offset_171; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6345 = _T_8 ? _GEN_1453 : offset_172; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6346 = _T_8 ? _GEN_1454 : offset_173; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6347 = _T_8 ? _GEN_1455 : offset_174; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6348 = _T_8 ? _GEN_1456 : offset_175; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6349 = _T_8 ? _GEN_1457 : offset_176; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6350 = _T_8 ? _GEN_1458 : offset_177; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6351 = _T_8 ? _GEN_1459 : offset_178; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6352 = _T_8 ? _GEN_1460 : offset_179; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6353 = _T_8 ? _GEN_1461 : offset_180; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6354 = _T_8 ? _GEN_1462 : offset_181; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6355 = _T_8 ? _GEN_1463 : offset_182; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6356 = _T_8 ? _GEN_1464 : offset_183; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6357 = _T_8 ? _GEN_1465 : offset_184; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6358 = _T_8 ? _GEN_1466 : offset_185; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6359 = _T_8 ? _GEN_1467 : offset_186; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6360 = _T_8 ? _GEN_1468 : offset_187; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6361 = _T_8 ? _GEN_1469 : offset_188; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6362 = _T_8 ? _GEN_1470 : offset_189; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6363 = _T_8 ? _GEN_1471 : offset_190; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6364 = _T_8 ? _GEN_1472 : offset_191; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6365 = _T_8 ? _GEN_1473 : offset_192; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6366 = _T_8 ? _GEN_1474 : offset_193; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6367 = _T_8 ? _GEN_1475 : offset_194; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6368 = _T_8 ? _GEN_1476 : offset_195; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6369 = _T_8 ? _GEN_1477 : offset_196; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6370 = _T_8 ? _GEN_1478 : offset_197; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6371 = _T_8 ? _GEN_1479 : offset_198; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6372 = _T_8 ? _GEN_1480 : offset_199; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6373 = _T_8 ? _GEN_1481 : offset_200; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6374 = _T_8 ? _GEN_1482 : offset_201; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6375 = _T_8 ? _GEN_1483 : offset_202; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6376 = _T_8 ? _GEN_1484 : offset_203; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6377 = _T_8 ? _GEN_1485 : offset_204; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6378 = _T_8 ? _GEN_1486 : offset_205; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6379 = _T_8 ? _GEN_1487 : offset_206; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6380 = _T_8 ? _GEN_1488 : offset_207; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6381 = _T_8 ? _GEN_1489 : offset_208; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6382 = _T_8 ? _GEN_1490 : offset_209; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6383 = _T_8 ? _GEN_1491 : offset_210; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6384 = _T_8 ? _GEN_1492 : offset_211; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6385 = _T_8 ? _GEN_1493 : offset_212; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6386 = _T_8 ? _GEN_1494 : offset_213; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6387 = _T_8 ? _GEN_1495 : offset_214; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6388 = _T_8 ? _GEN_1496 : offset_215; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6389 = _T_8 ? _GEN_1497 : offset_216; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6390 = _T_8 ? _GEN_1498 : offset_217; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6391 = _T_8 ? _GEN_1499 : offset_218; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6392 = _T_8 ? _GEN_1500 : offset_219; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6393 = _T_8 ? _GEN_1501 : offset_220; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6394 = _T_8 ? _GEN_1502 : offset_221; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6395 = _T_8 ? _GEN_1503 : offset_222; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6396 = _T_8 ? _GEN_1504 : offset_223; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6397 = _T_8 ? _GEN_1505 : offset_224; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6398 = _T_8 ? _GEN_1506 : offset_225; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6399 = _T_8 ? _GEN_1507 : offset_226; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6400 = _T_8 ? _GEN_1508 : offset_227; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6401 = _T_8 ? _GEN_1509 : offset_228; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6402 = _T_8 ? _GEN_1510 : offset_229; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6403 = _T_8 ? _GEN_1511 : offset_230; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6404 = _T_8 ? _GEN_1512 : offset_231; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6405 = _T_8 ? _GEN_1513 : offset_232; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6406 = _T_8 ? _GEN_1514 : offset_233; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6407 = _T_8 ? _GEN_1515 : offset_234; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6408 = _T_8 ? _GEN_1516 : offset_235; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6409 = _T_8 ? _GEN_1517 : offset_236; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6410 = _T_8 ? _GEN_1518 : offset_237; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6411 = _T_8 ? _GEN_1519 : offset_238; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6412 = _T_8 ? _GEN_1520 : offset_239; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6413 = _T_8 ? _GEN_1521 : offset_240; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6414 = _T_8 ? _GEN_1522 : offset_241; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6415 = _T_8 ? _GEN_1523 : offset_242; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6416 = _T_8 ? _GEN_1524 : offset_243; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6417 = _T_8 ? _GEN_1525 : offset_244; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6418 = _T_8 ? _GEN_1526 : offset_245; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6419 = _T_8 ? _GEN_1527 : offset_246; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6420 = _T_8 ? _GEN_1528 : offset_247; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6421 = _T_8 ? _GEN_1529 : offset_248; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6422 = _T_8 ? _GEN_1530 : offset_249; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6423 = _T_8 ? _GEN_1531 : offset_250; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6424 = _T_8 ? _GEN_1532 : offset_251; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6425 = _T_8 ? _GEN_1533 : offset_252; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6426 = _T_8 ? _GEN_1534 : offset_253; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6427 = _T_8 ? _GEN_1535 : offset_254; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6428 = _T_8 ? _GEN_1536 : offset_255; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [2:0] _GEN_6429 = _T_8 ? 3'h0 : state; // @[Conditional.scala 39:67 Dcache.scala 206:25 Dcache.scala 26:22]
  wire [2:0] _GEN_6430 = _T_6 ? _GEN_4366 : _GEN_6429; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_6431 = _T_6 ? _GEN_4367 : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_6437 = _T_6 ? _GEN_4373 : _GEN_5402; // @[Conditional.scala 39:67]
  wire  _GEN_6438 = _T_6 ? _GEN_4374 : _GEN_5404; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_6439 = _T_6 ? _GEN_4375 : cache_wdata; // @[Conditional.scala 39:67 Dcache.scala 118:28]
  wire [127:0] _GEN_6440 = _T_6 ? _GEN_4376 : cache_strb; // @[Conditional.scala 39:67 Dcache.scala 119:28]
  wire  _GEN_6441 = _T_6 ? data_ready : _GEN_5403; // @[Conditional.scala 39:67 Dcache.scala 46:28]
  wire  _GEN_6442 = _T_6 ? valid_0 : _GEN_5405; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6443 = _T_6 ? valid_1 : _GEN_5406; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6444 = _T_6 ? valid_2 : _GEN_5407; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6445 = _T_6 ? valid_3 : _GEN_5408; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6446 = _T_6 ? valid_4 : _GEN_5409; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6447 = _T_6 ? valid_5 : _GEN_5410; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6448 = _T_6 ? valid_6 : _GEN_5411; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6449 = _T_6 ? valid_7 : _GEN_5412; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6450 = _T_6 ? valid_8 : _GEN_5413; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6451 = _T_6 ? valid_9 : _GEN_5414; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6452 = _T_6 ? valid_10 : _GEN_5415; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6453 = _T_6 ? valid_11 : _GEN_5416; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6454 = _T_6 ? valid_12 : _GEN_5417; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6455 = _T_6 ? valid_13 : _GEN_5418; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6456 = _T_6 ? valid_14 : _GEN_5419; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6457 = _T_6 ? valid_15 : _GEN_5420; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6458 = _T_6 ? valid_16 : _GEN_5421; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6459 = _T_6 ? valid_17 : _GEN_5422; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6460 = _T_6 ? valid_18 : _GEN_5423; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6461 = _T_6 ? valid_19 : _GEN_5424; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6462 = _T_6 ? valid_20 : _GEN_5425; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6463 = _T_6 ? valid_21 : _GEN_5426; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6464 = _T_6 ? valid_22 : _GEN_5427; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6465 = _T_6 ? valid_23 : _GEN_5428; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6466 = _T_6 ? valid_24 : _GEN_5429; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6467 = _T_6 ? valid_25 : _GEN_5430; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6468 = _T_6 ? valid_26 : _GEN_5431; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6469 = _T_6 ? valid_27 : _GEN_5432; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6470 = _T_6 ? valid_28 : _GEN_5433; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6471 = _T_6 ? valid_29 : _GEN_5434; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6472 = _T_6 ? valid_30 : _GEN_5435; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6473 = _T_6 ? valid_31 : _GEN_5436; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6474 = _T_6 ? valid_32 : _GEN_5437; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6475 = _T_6 ? valid_33 : _GEN_5438; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6476 = _T_6 ? valid_34 : _GEN_5439; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6477 = _T_6 ? valid_35 : _GEN_5440; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6478 = _T_6 ? valid_36 : _GEN_5441; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6479 = _T_6 ? valid_37 : _GEN_5442; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6480 = _T_6 ? valid_38 : _GEN_5443; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6481 = _T_6 ? valid_39 : _GEN_5444; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6482 = _T_6 ? valid_40 : _GEN_5445; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6483 = _T_6 ? valid_41 : _GEN_5446; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6484 = _T_6 ? valid_42 : _GEN_5447; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6485 = _T_6 ? valid_43 : _GEN_5448; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6486 = _T_6 ? valid_44 : _GEN_5449; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6487 = _T_6 ? valid_45 : _GEN_5450; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6488 = _T_6 ? valid_46 : _GEN_5451; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6489 = _T_6 ? valid_47 : _GEN_5452; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6490 = _T_6 ? valid_48 : _GEN_5453; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6491 = _T_6 ? valid_49 : _GEN_5454; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6492 = _T_6 ? valid_50 : _GEN_5455; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6493 = _T_6 ? valid_51 : _GEN_5456; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6494 = _T_6 ? valid_52 : _GEN_5457; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6495 = _T_6 ? valid_53 : _GEN_5458; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6496 = _T_6 ? valid_54 : _GEN_5459; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6497 = _T_6 ? valid_55 : _GEN_5460; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6498 = _T_6 ? valid_56 : _GEN_5461; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6499 = _T_6 ? valid_57 : _GEN_5462; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6500 = _T_6 ? valid_58 : _GEN_5463; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6501 = _T_6 ? valid_59 : _GEN_5464; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6502 = _T_6 ? valid_60 : _GEN_5465; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6503 = _T_6 ? valid_61 : _GEN_5466; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6504 = _T_6 ? valid_62 : _GEN_5467; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6505 = _T_6 ? valid_63 : _GEN_5468; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6506 = _T_6 ? valid_64 : _GEN_5469; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6507 = _T_6 ? valid_65 : _GEN_5470; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6508 = _T_6 ? valid_66 : _GEN_5471; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6509 = _T_6 ? valid_67 : _GEN_5472; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6510 = _T_6 ? valid_68 : _GEN_5473; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6511 = _T_6 ? valid_69 : _GEN_5474; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6512 = _T_6 ? valid_70 : _GEN_5475; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6513 = _T_6 ? valid_71 : _GEN_5476; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6514 = _T_6 ? valid_72 : _GEN_5477; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6515 = _T_6 ? valid_73 : _GEN_5478; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6516 = _T_6 ? valid_74 : _GEN_5479; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6517 = _T_6 ? valid_75 : _GEN_5480; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6518 = _T_6 ? valid_76 : _GEN_5481; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6519 = _T_6 ? valid_77 : _GEN_5482; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6520 = _T_6 ? valid_78 : _GEN_5483; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6521 = _T_6 ? valid_79 : _GEN_5484; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6522 = _T_6 ? valid_80 : _GEN_5485; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6523 = _T_6 ? valid_81 : _GEN_5486; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6524 = _T_6 ? valid_82 : _GEN_5487; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6525 = _T_6 ? valid_83 : _GEN_5488; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6526 = _T_6 ? valid_84 : _GEN_5489; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6527 = _T_6 ? valid_85 : _GEN_5490; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6528 = _T_6 ? valid_86 : _GEN_5491; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6529 = _T_6 ? valid_87 : _GEN_5492; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6530 = _T_6 ? valid_88 : _GEN_5493; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6531 = _T_6 ? valid_89 : _GEN_5494; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6532 = _T_6 ? valid_90 : _GEN_5495; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6533 = _T_6 ? valid_91 : _GEN_5496; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6534 = _T_6 ? valid_92 : _GEN_5497; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6535 = _T_6 ? valid_93 : _GEN_5498; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6536 = _T_6 ? valid_94 : _GEN_5499; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6537 = _T_6 ? valid_95 : _GEN_5500; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6538 = _T_6 ? valid_96 : _GEN_5501; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6539 = _T_6 ? valid_97 : _GEN_5502; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6540 = _T_6 ? valid_98 : _GEN_5503; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6541 = _T_6 ? valid_99 : _GEN_5504; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6542 = _T_6 ? valid_100 : _GEN_5505; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6543 = _T_6 ? valid_101 : _GEN_5506; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6544 = _T_6 ? valid_102 : _GEN_5507; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6545 = _T_6 ? valid_103 : _GEN_5508; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6546 = _T_6 ? valid_104 : _GEN_5509; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6547 = _T_6 ? valid_105 : _GEN_5510; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6548 = _T_6 ? valid_106 : _GEN_5511; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6549 = _T_6 ? valid_107 : _GEN_5512; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6550 = _T_6 ? valid_108 : _GEN_5513; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6551 = _T_6 ? valid_109 : _GEN_5514; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6552 = _T_6 ? valid_110 : _GEN_5515; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6553 = _T_6 ? valid_111 : _GEN_5516; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6554 = _T_6 ? valid_112 : _GEN_5517; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6555 = _T_6 ? valid_113 : _GEN_5518; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6556 = _T_6 ? valid_114 : _GEN_5519; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6557 = _T_6 ? valid_115 : _GEN_5520; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6558 = _T_6 ? valid_116 : _GEN_5521; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6559 = _T_6 ? valid_117 : _GEN_5522; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6560 = _T_6 ? valid_118 : _GEN_5523; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6561 = _T_6 ? valid_119 : _GEN_5524; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6562 = _T_6 ? valid_120 : _GEN_5525; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6563 = _T_6 ? valid_121 : _GEN_5526; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6564 = _T_6 ? valid_122 : _GEN_5527; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6565 = _T_6 ? valid_123 : _GEN_5528; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6566 = _T_6 ? valid_124 : _GEN_5529; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6567 = _T_6 ? valid_125 : _GEN_5530; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6568 = _T_6 ? valid_126 : _GEN_5531; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6569 = _T_6 ? valid_127 : _GEN_5532; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6570 = _T_6 ? valid_128 : _GEN_5533; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6571 = _T_6 ? valid_129 : _GEN_5534; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6572 = _T_6 ? valid_130 : _GEN_5535; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6573 = _T_6 ? valid_131 : _GEN_5536; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6574 = _T_6 ? valid_132 : _GEN_5537; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6575 = _T_6 ? valid_133 : _GEN_5538; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6576 = _T_6 ? valid_134 : _GEN_5539; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6577 = _T_6 ? valid_135 : _GEN_5540; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6578 = _T_6 ? valid_136 : _GEN_5541; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6579 = _T_6 ? valid_137 : _GEN_5542; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6580 = _T_6 ? valid_138 : _GEN_5543; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6581 = _T_6 ? valid_139 : _GEN_5544; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6582 = _T_6 ? valid_140 : _GEN_5545; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6583 = _T_6 ? valid_141 : _GEN_5546; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6584 = _T_6 ? valid_142 : _GEN_5547; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6585 = _T_6 ? valid_143 : _GEN_5548; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6586 = _T_6 ? valid_144 : _GEN_5549; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6587 = _T_6 ? valid_145 : _GEN_5550; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6588 = _T_6 ? valid_146 : _GEN_5551; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6589 = _T_6 ? valid_147 : _GEN_5552; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6590 = _T_6 ? valid_148 : _GEN_5553; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6591 = _T_6 ? valid_149 : _GEN_5554; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6592 = _T_6 ? valid_150 : _GEN_5555; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6593 = _T_6 ? valid_151 : _GEN_5556; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6594 = _T_6 ? valid_152 : _GEN_5557; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6595 = _T_6 ? valid_153 : _GEN_5558; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6596 = _T_6 ? valid_154 : _GEN_5559; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6597 = _T_6 ? valid_155 : _GEN_5560; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6598 = _T_6 ? valid_156 : _GEN_5561; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6599 = _T_6 ? valid_157 : _GEN_5562; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6600 = _T_6 ? valid_158 : _GEN_5563; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6601 = _T_6 ? valid_159 : _GEN_5564; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6602 = _T_6 ? valid_160 : _GEN_5565; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6603 = _T_6 ? valid_161 : _GEN_5566; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6604 = _T_6 ? valid_162 : _GEN_5567; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6605 = _T_6 ? valid_163 : _GEN_5568; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6606 = _T_6 ? valid_164 : _GEN_5569; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6607 = _T_6 ? valid_165 : _GEN_5570; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6608 = _T_6 ? valid_166 : _GEN_5571; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6609 = _T_6 ? valid_167 : _GEN_5572; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6610 = _T_6 ? valid_168 : _GEN_5573; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6611 = _T_6 ? valid_169 : _GEN_5574; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6612 = _T_6 ? valid_170 : _GEN_5575; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6613 = _T_6 ? valid_171 : _GEN_5576; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6614 = _T_6 ? valid_172 : _GEN_5577; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6615 = _T_6 ? valid_173 : _GEN_5578; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6616 = _T_6 ? valid_174 : _GEN_5579; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6617 = _T_6 ? valid_175 : _GEN_5580; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6618 = _T_6 ? valid_176 : _GEN_5581; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6619 = _T_6 ? valid_177 : _GEN_5582; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6620 = _T_6 ? valid_178 : _GEN_5583; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6621 = _T_6 ? valid_179 : _GEN_5584; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6622 = _T_6 ? valid_180 : _GEN_5585; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6623 = _T_6 ? valid_181 : _GEN_5586; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6624 = _T_6 ? valid_182 : _GEN_5587; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6625 = _T_6 ? valid_183 : _GEN_5588; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6626 = _T_6 ? valid_184 : _GEN_5589; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6627 = _T_6 ? valid_185 : _GEN_5590; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6628 = _T_6 ? valid_186 : _GEN_5591; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6629 = _T_6 ? valid_187 : _GEN_5592; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6630 = _T_6 ? valid_188 : _GEN_5593; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6631 = _T_6 ? valid_189 : _GEN_5594; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6632 = _T_6 ? valid_190 : _GEN_5595; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6633 = _T_6 ? valid_191 : _GEN_5596; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6634 = _T_6 ? valid_192 : _GEN_5597; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6635 = _T_6 ? valid_193 : _GEN_5598; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6636 = _T_6 ? valid_194 : _GEN_5599; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6637 = _T_6 ? valid_195 : _GEN_5600; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6638 = _T_6 ? valid_196 : _GEN_5601; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6639 = _T_6 ? valid_197 : _GEN_5602; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6640 = _T_6 ? valid_198 : _GEN_5603; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6641 = _T_6 ? valid_199 : _GEN_5604; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6642 = _T_6 ? valid_200 : _GEN_5605; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6643 = _T_6 ? valid_201 : _GEN_5606; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6644 = _T_6 ? valid_202 : _GEN_5607; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6645 = _T_6 ? valid_203 : _GEN_5608; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6646 = _T_6 ? valid_204 : _GEN_5609; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6647 = _T_6 ? valid_205 : _GEN_5610; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6648 = _T_6 ? valid_206 : _GEN_5611; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6649 = _T_6 ? valid_207 : _GEN_5612; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6650 = _T_6 ? valid_208 : _GEN_5613; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6651 = _T_6 ? valid_209 : _GEN_5614; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6652 = _T_6 ? valid_210 : _GEN_5615; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6653 = _T_6 ? valid_211 : _GEN_5616; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6654 = _T_6 ? valid_212 : _GEN_5617; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6655 = _T_6 ? valid_213 : _GEN_5618; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6656 = _T_6 ? valid_214 : _GEN_5619; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6657 = _T_6 ? valid_215 : _GEN_5620; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6658 = _T_6 ? valid_216 : _GEN_5621; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6659 = _T_6 ? valid_217 : _GEN_5622; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6660 = _T_6 ? valid_218 : _GEN_5623; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6661 = _T_6 ? valid_219 : _GEN_5624; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6662 = _T_6 ? valid_220 : _GEN_5625; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6663 = _T_6 ? valid_221 : _GEN_5626; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6664 = _T_6 ? valid_222 : _GEN_5627; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6665 = _T_6 ? valid_223 : _GEN_5628; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6666 = _T_6 ? valid_224 : _GEN_5629; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6667 = _T_6 ? valid_225 : _GEN_5630; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6668 = _T_6 ? valid_226 : _GEN_5631; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6669 = _T_6 ? valid_227 : _GEN_5632; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6670 = _T_6 ? valid_228 : _GEN_5633; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6671 = _T_6 ? valid_229 : _GEN_5634; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6672 = _T_6 ? valid_230 : _GEN_5635; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6673 = _T_6 ? valid_231 : _GEN_5636; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6674 = _T_6 ? valid_232 : _GEN_5637; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6675 = _T_6 ? valid_233 : _GEN_5638; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6676 = _T_6 ? valid_234 : _GEN_5639; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6677 = _T_6 ? valid_235 : _GEN_5640; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6678 = _T_6 ? valid_236 : _GEN_5641; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6679 = _T_6 ? valid_237 : _GEN_5642; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6680 = _T_6 ? valid_238 : _GEN_5643; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6681 = _T_6 ? valid_239 : _GEN_5644; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6682 = _T_6 ? valid_240 : _GEN_5645; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6683 = _T_6 ? valid_241 : _GEN_5646; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6684 = _T_6 ? valid_242 : _GEN_5647; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6685 = _T_6 ? valid_243 : _GEN_5648; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6686 = _T_6 ? valid_244 : _GEN_5649; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6687 = _T_6 ? valid_245 : _GEN_5650; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6688 = _T_6 ? valid_246 : _GEN_5651; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6689 = _T_6 ? valid_247 : _GEN_5652; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6690 = _T_6 ? valid_248 : _GEN_5653; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6691 = _T_6 ? valid_249 : _GEN_5654; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6692 = _T_6 ? valid_250 : _GEN_5655; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6693 = _T_6 ? valid_251 : _GEN_5656; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6694 = _T_6 ? valid_252 : _GEN_5657; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6695 = _T_6 ? valid_253 : _GEN_5658; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6696 = _T_6 ? valid_254 : _GEN_5659; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6697 = _T_6 ? valid_255 : _GEN_5660; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire [19:0] _GEN_6698 = _T_6 ? tag_0 : _GEN_5661; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6699 = _T_6 ? tag_1 : _GEN_5662; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6700 = _T_6 ? tag_2 : _GEN_5663; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6701 = _T_6 ? tag_3 : _GEN_5664; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6702 = _T_6 ? tag_4 : _GEN_5665; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6703 = _T_6 ? tag_5 : _GEN_5666; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6704 = _T_6 ? tag_6 : _GEN_5667; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6705 = _T_6 ? tag_7 : _GEN_5668; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6706 = _T_6 ? tag_8 : _GEN_5669; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6707 = _T_6 ? tag_9 : _GEN_5670; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6708 = _T_6 ? tag_10 : _GEN_5671; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6709 = _T_6 ? tag_11 : _GEN_5672; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6710 = _T_6 ? tag_12 : _GEN_5673; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6711 = _T_6 ? tag_13 : _GEN_5674; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6712 = _T_6 ? tag_14 : _GEN_5675; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6713 = _T_6 ? tag_15 : _GEN_5676; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6714 = _T_6 ? tag_16 : _GEN_5677; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6715 = _T_6 ? tag_17 : _GEN_5678; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6716 = _T_6 ? tag_18 : _GEN_5679; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6717 = _T_6 ? tag_19 : _GEN_5680; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6718 = _T_6 ? tag_20 : _GEN_5681; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6719 = _T_6 ? tag_21 : _GEN_5682; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6720 = _T_6 ? tag_22 : _GEN_5683; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6721 = _T_6 ? tag_23 : _GEN_5684; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6722 = _T_6 ? tag_24 : _GEN_5685; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6723 = _T_6 ? tag_25 : _GEN_5686; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6724 = _T_6 ? tag_26 : _GEN_5687; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6725 = _T_6 ? tag_27 : _GEN_5688; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6726 = _T_6 ? tag_28 : _GEN_5689; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6727 = _T_6 ? tag_29 : _GEN_5690; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6728 = _T_6 ? tag_30 : _GEN_5691; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6729 = _T_6 ? tag_31 : _GEN_5692; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6730 = _T_6 ? tag_32 : _GEN_5693; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6731 = _T_6 ? tag_33 : _GEN_5694; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6732 = _T_6 ? tag_34 : _GEN_5695; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6733 = _T_6 ? tag_35 : _GEN_5696; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6734 = _T_6 ? tag_36 : _GEN_5697; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6735 = _T_6 ? tag_37 : _GEN_5698; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6736 = _T_6 ? tag_38 : _GEN_5699; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6737 = _T_6 ? tag_39 : _GEN_5700; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6738 = _T_6 ? tag_40 : _GEN_5701; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6739 = _T_6 ? tag_41 : _GEN_5702; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6740 = _T_6 ? tag_42 : _GEN_5703; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6741 = _T_6 ? tag_43 : _GEN_5704; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6742 = _T_6 ? tag_44 : _GEN_5705; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6743 = _T_6 ? tag_45 : _GEN_5706; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6744 = _T_6 ? tag_46 : _GEN_5707; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6745 = _T_6 ? tag_47 : _GEN_5708; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6746 = _T_6 ? tag_48 : _GEN_5709; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6747 = _T_6 ? tag_49 : _GEN_5710; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6748 = _T_6 ? tag_50 : _GEN_5711; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6749 = _T_6 ? tag_51 : _GEN_5712; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6750 = _T_6 ? tag_52 : _GEN_5713; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6751 = _T_6 ? tag_53 : _GEN_5714; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6752 = _T_6 ? tag_54 : _GEN_5715; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6753 = _T_6 ? tag_55 : _GEN_5716; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6754 = _T_6 ? tag_56 : _GEN_5717; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6755 = _T_6 ? tag_57 : _GEN_5718; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6756 = _T_6 ? tag_58 : _GEN_5719; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6757 = _T_6 ? tag_59 : _GEN_5720; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6758 = _T_6 ? tag_60 : _GEN_5721; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6759 = _T_6 ? tag_61 : _GEN_5722; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6760 = _T_6 ? tag_62 : _GEN_5723; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6761 = _T_6 ? tag_63 : _GEN_5724; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6762 = _T_6 ? tag_64 : _GEN_5725; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6763 = _T_6 ? tag_65 : _GEN_5726; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6764 = _T_6 ? tag_66 : _GEN_5727; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6765 = _T_6 ? tag_67 : _GEN_5728; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6766 = _T_6 ? tag_68 : _GEN_5729; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6767 = _T_6 ? tag_69 : _GEN_5730; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6768 = _T_6 ? tag_70 : _GEN_5731; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6769 = _T_6 ? tag_71 : _GEN_5732; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6770 = _T_6 ? tag_72 : _GEN_5733; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6771 = _T_6 ? tag_73 : _GEN_5734; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6772 = _T_6 ? tag_74 : _GEN_5735; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6773 = _T_6 ? tag_75 : _GEN_5736; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6774 = _T_6 ? tag_76 : _GEN_5737; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6775 = _T_6 ? tag_77 : _GEN_5738; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6776 = _T_6 ? tag_78 : _GEN_5739; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6777 = _T_6 ? tag_79 : _GEN_5740; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6778 = _T_6 ? tag_80 : _GEN_5741; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6779 = _T_6 ? tag_81 : _GEN_5742; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6780 = _T_6 ? tag_82 : _GEN_5743; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6781 = _T_6 ? tag_83 : _GEN_5744; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6782 = _T_6 ? tag_84 : _GEN_5745; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6783 = _T_6 ? tag_85 : _GEN_5746; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6784 = _T_6 ? tag_86 : _GEN_5747; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6785 = _T_6 ? tag_87 : _GEN_5748; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6786 = _T_6 ? tag_88 : _GEN_5749; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6787 = _T_6 ? tag_89 : _GEN_5750; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6788 = _T_6 ? tag_90 : _GEN_5751; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6789 = _T_6 ? tag_91 : _GEN_5752; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6790 = _T_6 ? tag_92 : _GEN_5753; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6791 = _T_6 ? tag_93 : _GEN_5754; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6792 = _T_6 ? tag_94 : _GEN_5755; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6793 = _T_6 ? tag_95 : _GEN_5756; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6794 = _T_6 ? tag_96 : _GEN_5757; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6795 = _T_6 ? tag_97 : _GEN_5758; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6796 = _T_6 ? tag_98 : _GEN_5759; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6797 = _T_6 ? tag_99 : _GEN_5760; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6798 = _T_6 ? tag_100 : _GEN_5761; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6799 = _T_6 ? tag_101 : _GEN_5762; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6800 = _T_6 ? tag_102 : _GEN_5763; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6801 = _T_6 ? tag_103 : _GEN_5764; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6802 = _T_6 ? tag_104 : _GEN_5765; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6803 = _T_6 ? tag_105 : _GEN_5766; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6804 = _T_6 ? tag_106 : _GEN_5767; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6805 = _T_6 ? tag_107 : _GEN_5768; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6806 = _T_6 ? tag_108 : _GEN_5769; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6807 = _T_6 ? tag_109 : _GEN_5770; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6808 = _T_6 ? tag_110 : _GEN_5771; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6809 = _T_6 ? tag_111 : _GEN_5772; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6810 = _T_6 ? tag_112 : _GEN_5773; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6811 = _T_6 ? tag_113 : _GEN_5774; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6812 = _T_6 ? tag_114 : _GEN_5775; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6813 = _T_6 ? tag_115 : _GEN_5776; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6814 = _T_6 ? tag_116 : _GEN_5777; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6815 = _T_6 ? tag_117 : _GEN_5778; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6816 = _T_6 ? tag_118 : _GEN_5779; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6817 = _T_6 ? tag_119 : _GEN_5780; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6818 = _T_6 ? tag_120 : _GEN_5781; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6819 = _T_6 ? tag_121 : _GEN_5782; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6820 = _T_6 ? tag_122 : _GEN_5783; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6821 = _T_6 ? tag_123 : _GEN_5784; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6822 = _T_6 ? tag_124 : _GEN_5785; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6823 = _T_6 ? tag_125 : _GEN_5786; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6824 = _T_6 ? tag_126 : _GEN_5787; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6825 = _T_6 ? tag_127 : _GEN_5788; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6826 = _T_6 ? tag_128 : _GEN_5789; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6827 = _T_6 ? tag_129 : _GEN_5790; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6828 = _T_6 ? tag_130 : _GEN_5791; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6829 = _T_6 ? tag_131 : _GEN_5792; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6830 = _T_6 ? tag_132 : _GEN_5793; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6831 = _T_6 ? tag_133 : _GEN_5794; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6832 = _T_6 ? tag_134 : _GEN_5795; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6833 = _T_6 ? tag_135 : _GEN_5796; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6834 = _T_6 ? tag_136 : _GEN_5797; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6835 = _T_6 ? tag_137 : _GEN_5798; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6836 = _T_6 ? tag_138 : _GEN_5799; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6837 = _T_6 ? tag_139 : _GEN_5800; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6838 = _T_6 ? tag_140 : _GEN_5801; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6839 = _T_6 ? tag_141 : _GEN_5802; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6840 = _T_6 ? tag_142 : _GEN_5803; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6841 = _T_6 ? tag_143 : _GEN_5804; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6842 = _T_6 ? tag_144 : _GEN_5805; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6843 = _T_6 ? tag_145 : _GEN_5806; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6844 = _T_6 ? tag_146 : _GEN_5807; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6845 = _T_6 ? tag_147 : _GEN_5808; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6846 = _T_6 ? tag_148 : _GEN_5809; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6847 = _T_6 ? tag_149 : _GEN_5810; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6848 = _T_6 ? tag_150 : _GEN_5811; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6849 = _T_6 ? tag_151 : _GEN_5812; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6850 = _T_6 ? tag_152 : _GEN_5813; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6851 = _T_6 ? tag_153 : _GEN_5814; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6852 = _T_6 ? tag_154 : _GEN_5815; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6853 = _T_6 ? tag_155 : _GEN_5816; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6854 = _T_6 ? tag_156 : _GEN_5817; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6855 = _T_6 ? tag_157 : _GEN_5818; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6856 = _T_6 ? tag_158 : _GEN_5819; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6857 = _T_6 ? tag_159 : _GEN_5820; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6858 = _T_6 ? tag_160 : _GEN_5821; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6859 = _T_6 ? tag_161 : _GEN_5822; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6860 = _T_6 ? tag_162 : _GEN_5823; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6861 = _T_6 ? tag_163 : _GEN_5824; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6862 = _T_6 ? tag_164 : _GEN_5825; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6863 = _T_6 ? tag_165 : _GEN_5826; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6864 = _T_6 ? tag_166 : _GEN_5827; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6865 = _T_6 ? tag_167 : _GEN_5828; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6866 = _T_6 ? tag_168 : _GEN_5829; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6867 = _T_6 ? tag_169 : _GEN_5830; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6868 = _T_6 ? tag_170 : _GEN_5831; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6869 = _T_6 ? tag_171 : _GEN_5832; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6870 = _T_6 ? tag_172 : _GEN_5833; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6871 = _T_6 ? tag_173 : _GEN_5834; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6872 = _T_6 ? tag_174 : _GEN_5835; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6873 = _T_6 ? tag_175 : _GEN_5836; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6874 = _T_6 ? tag_176 : _GEN_5837; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6875 = _T_6 ? tag_177 : _GEN_5838; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6876 = _T_6 ? tag_178 : _GEN_5839; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6877 = _T_6 ? tag_179 : _GEN_5840; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6878 = _T_6 ? tag_180 : _GEN_5841; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6879 = _T_6 ? tag_181 : _GEN_5842; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6880 = _T_6 ? tag_182 : _GEN_5843; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6881 = _T_6 ? tag_183 : _GEN_5844; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6882 = _T_6 ? tag_184 : _GEN_5845; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6883 = _T_6 ? tag_185 : _GEN_5846; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6884 = _T_6 ? tag_186 : _GEN_5847; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6885 = _T_6 ? tag_187 : _GEN_5848; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6886 = _T_6 ? tag_188 : _GEN_5849; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6887 = _T_6 ? tag_189 : _GEN_5850; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6888 = _T_6 ? tag_190 : _GEN_5851; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6889 = _T_6 ? tag_191 : _GEN_5852; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6890 = _T_6 ? tag_192 : _GEN_5853; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6891 = _T_6 ? tag_193 : _GEN_5854; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6892 = _T_6 ? tag_194 : _GEN_5855; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6893 = _T_6 ? tag_195 : _GEN_5856; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6894 = _T_6 ? tag_196 : _GEN_5857; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6895 = _T_6 ? tag_197 : _GEN_5858; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6896 = _T_6 ? tag_198 : _GEN_5859; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6897 = _T_6 ? tag_199 : _GEN_5860; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6898 = _T_6 ? tag_200 : _GEN_5861; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6899 = _T_6 ? tag_201 : _GEN_5862; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6900 = _T_6 ? tag_202 : _GEN_5863; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6901 = _T_6 ? tag_203 : _GEN_5864; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6902 = _T_6 ? tag_204 : _GEN_5865; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6903 = _T_6 ? tag_205 : _GEN_5866; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6904 = _T_6 ? tag_206 : _GEN_5867; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6905 = _T_6 ? tag_207 : _GEN_5868; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6906 = _T_6 ? tag_208 : _GEN_5869; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6907 = _T_6 ? tag_209 : _GEN_5870; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6908 = _T_6 ? tag_210 : _GEN_5871; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6909 = _T_6 ? tag_211 : _GEN_5872; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6910 = _T_6 ? tag_212 : _GEN_5873; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6911 = _T_6 ? tag_213 : _GEN_5874; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6912 = _T_6 ? tag_214 : _GEN_5875; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6913 = _T_6 ? tag_215 : _GEN_5876; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6914 = _T_6 ? tag_216 : _GEN_5877; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6915 = _T_6 ? tag_217 : _GEN_5878; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6916 = _T_6 ? tag_218 : _GEN_5879; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6917 = _T_6 ? tag_219 : _GEN_5880; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6918 = _T_6 ? tag_220 : _GEN_5881; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6919 = _T_6 ? tag_221 : _GEN_5882; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6920 = _T_6 ? tag_222 : _GEN_5883; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6921 = _T_6 ? tag_223 : _GEN_5884; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6922 = _T_6 ? tag_224 : _GEN_5885; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6923 = _T_6 ? tag_225 : _GEN_5886; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6924 = _T_6 ? tag_226 : _GEN_5887; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6925 = _T_6 ? tag_227 : _GEN_5888; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6926 = _T_6 ? tag_228 : _GEN_5889; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6927 = _T_6 ? tag_229 : _GEN_5890; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6928 = _T_6 ? tag_230 : _GEN_5891; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6929 = _T_6 ? tag_231 : _GEN_5892; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6930 = _T_6 ? tag_232 : _GEN_5893; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6931 = _T_6 ? tag_233 : _GEN_5894; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6932 = _T_6 ? tag_234 : _GEN_5895; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6933 = _T_6 ? tag_235 : _GEN_5896; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6934 = _T_6 ? tag_236 : _GEN_5897; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6935 = _T_6 ? tag_237 : _GEN_5898; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6936 = _T_6 ? tag_238 : _GEN_5899; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6937 = _T_6 ? tag_239 : _GEN_5900; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6938 = _T_6 ? tag_240 : _GEN_5901; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6939 = _T_6 ? tag_241 : _GEN_5902; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6940 = _T_6 ? tag_242 : _GEN_5903; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6941 = _T_6 ? tag_243 : _GEN_5904; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6942 = _T_6 ? tag_244 : _GEN_5905; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6943 = _T_6 ? tag_245 : _GEN_5906; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6944 = _T_6 ? tag_246 : _GEN_5907; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6945 = _T_6 ? tag_247 : _GEN_5908; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6946 = _T_6 ? tag_248 : _GEN_5909; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6947 = _T_6 ? tag_249 : _GEN_5910; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6948 = _T_6 ? tag_250 : _GEN_5911; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6949 = _T_6 ? tag_251 : _GEN_5912; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6950 = _T_6 ? tag_252 : _GEN_5913; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6951 = _T_6 ? tag_253 : _GEN_5914; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6952 = _T_6 ? tag_254 : _GEN_5915; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6953 = _T_6 ? tag_255 : _GEN_5916; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire  _GEN_6954 = _T_6 ? dirty_0 : _GEN_5917; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6955 = _T_6 ? dirty_1 : _GEN_5918; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6956 = _T_6 ? dirty_2 : _GEN_5919; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6957 = _T_6 ? dirty_3 : _GEN_5920; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6958 = _T_6 ? dirty_4 : _GEN_5921; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6959 = _T_6 ? dirty_5 : _GEN_5922; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6960 = _T_6 ? dirty_6 : _GEN_5923; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6961 = _T_6 ? dirty_7 : _GEN_5924; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6962 = _T_6 ? dirty_8 : _GEN_5925; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6963 = _T_6 ? dirty_9 : _GEN_5926; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6964 = _T_6 ? dirty_10 : _GEN_5927; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6965 = _T_6 ? dirty_11 : _GEN_5928; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6966 = _T_6 ? dirty_12 : _GEN_5929; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6967 = _T_6 ? dirty_13 : _GEN_5930; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6968 = _T_6 ? dirty_14 : _GEN_5931; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6969 = _T_6 ? dirty_15 : _GEN_5932; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6970 = _T_6 ? dirty_16 : _GEN_5933; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6971 = _T_6 ? dirty_17 : _GEN_5934; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6972 = _T_6 ? dirty_18 : _GEN_5935; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6973 = _T_6 ? dirty_19 : _GEN_5936; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6974 = _T_6 ? dirty_20 : _GEN_5937; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6975 = _T_6 ? dirty_21 : _GEN_5938; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6976 = _T_6 ? dirty_22 : _GEN_5939; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6977 = _T_6 ? dirty_23 : _GEN_5940; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6978 = _T_6 ? dirty_24 : _GEN_5941; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6979 = _T_6 ? dirty_25 : _GEN_5942; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6980 = _T_6 ? dirty_26 : _GEN_5943; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6981 = _T_6 ? dirty_27 : _GEN_5944; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6982 = _T_6 ? dirty_28 : _GEN_5945; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6983 = _T_6 ? dirty_29 : _GEN_5946; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6984 = _T_6 ? dirty_30 : _GEN_5947; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6985 = _T_6 ? dirty_31 : _GEN_5948; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6986 = _T_6 ? dirty_32 : _GEN_5949; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6987 = _T_6 ? dirty_33 : _GEN_5950; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6988 = _T_6 ? dirty_34 : _GEN_5951; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6989 = _T_6 ? dirty_35 : _GEN_5952; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6990 = _T_6 ? dirty_36 : _GEN_5953; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6991 = _T_6 ? dirty_37 : _GEN_5954; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6992 = _T_6 ? dirty_38 : _GEN_5955; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6993 = _T_6 ? dirty_39 : _GEN_5956; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6994 = _T_6 ? dirty_40 : _GEN_5957; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6995 = _T_6 ? dirty_41 : _GEN_5958; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6996 = _T_6 ? dirty_42 : _GEN_5959; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6997 = _T_6 ? dirty_43 : _GEN_5960; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6998 = _T_6 ? dirty_44 : _GEN_5961; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6999 = _T_6 ? dirty_45 : _GEN_5962; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7000 = _T_6 ? dirty_46 : _GEN_5963; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7001 = _T_6 ? dirty_47 : _GEN_5964; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7002 = _T_6 ? dirty_48 : _GEN_5965; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7003 = _T_6 ? dirty_49 : _GEN_5966; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7004 = _T_6 ? dirty_50 : _GEN_5967; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7005 = _T_6 ? dirty_51 : _GEN_5968; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7006 = _T_6 ? dirty_52 : _GEN_5969; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7007 = _T_6 ? dirty_53 : _GEN_5970; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7008 = _T_6 ? dirty_54 : _GEN_5971; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7009 = _T_6 ? dirty_55 : _GEN_5972; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7010 = _T_6 ? dirty_56 : _GEN_5973; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7011 = _T_6 ? dirty_57 : _GEN_5974; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7012 = _T_6 ? dirty_58 : _GEN_5975; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7013 = _T_6 ? dirty_59 : _GEN_5976; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7014 = _T_6 ? dirty_60 : _GEN_5977; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7015 = _T_6 ? dirty_61 : _GEN_5978; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7016 = _T_6 ? dirty_62 : _GEN_5979; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7017 = _T_6 ? dirty_63 : _GEN_5980; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7018 = _T_6 ? dirty_64 : _GEN_5981; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7019 = _T_6 ? dirty_65 : _GEN_5982; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7020 = _T_6 ? dirty_66 : _GEN_5983; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7021 = _T_6 ? dirty_67 : _GEN_5984; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7022 = _T_6 ? dirty_68 : _GEN_5985; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7023 = _T_6 ? dirty_69 : _GEN_5986; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7024 = _T_6 ? dirty_70 : _GEN_5987; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7025 = _T_6 ? dirty_71 : _GEN_5988; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7026 = _T_6 ? dirty_72 : _GEN_5989; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7027 = _T_6 ? dirty_73 : _GEN_5990; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7028 = _T_6 ? dirty_74 : _GEN_5991; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7029 = _T_6 ? dirty_75 : _GEN_5992; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7030 = _T_6 ? dirty_76 : _GEN_5993; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7031 = _T_6 ? dirty_77 : _GEN_5994; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7032 = _T_6 ? dirty_78 : _GEN_5995; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7033 = _T_6 ? dirty_79 : _GEN_5996; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7034 = _T_6 ? dirty_80 : _GEN_5997; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7035 = _T_6 ? dirty_81 : _GEN_5998; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7036 = _T_6 ? dirty_82 : _GEN_5999; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7037 = _T_6 ? dirty_83 : _GEN_6000; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7038 = _T_6 ? dirty_84 : _GEN_6001; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7039 = _T_6 ? dirty_85 : _GEN_6002; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7040 = _T_6 ? dirty_86 : _GEN_6003; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7041 = _T_6 ? dirty_87 : _GEN_6004; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7042 = _T_6 ? dirty_88 : _GEN_6005; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7043 = _T_6 ? dirty_89 : _GEN_6006; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7044 = _T_6 ? dirty_90 : _GEN_6007; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7045 = _T_6 ? dirty_91 : _GEN_6008; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7046 = _T_6 ? dirty_92 : _GEN_6009; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7047 = _T_6 ? dirty_93 : _GEN_6010; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7048 = _T_6 ? dirty_94 : _GEN_6011; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7049 = _T_6 ? dirty_95 : _GEN_6012; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7050 = _T_6 ? dirty_96 : _GEN_6013; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7051 = _T_6 ? dirty_97 : _GEN_6014; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7052 = _T_6 ? dirty_98 : _GEN_6015; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7053 = _T_6 ? dirty_99 : _GEN_6016; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7054 = _T_6 ? dirty_100 : _GEN_6017; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7055 = _T_6 ? dirty_101 : _GEN_6018; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7056 = _T_6 ? dirty_102 : _GEN_6019; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7057 = _T_6 ? dirty_103 : _GEN_6020; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7058 = _T_6 ? dirty_104 : _GEN_6021; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7059 = _T_6 ? dirty_105 : _GEN_6022; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7060 = _T_6 ? dirty_106 : _GEN_6023; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7061 = _T_6 ? dirty_107 : _GEN_6024; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7062 = _T_6 ? dirty_108 : _GEN_6025; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7063 = _T_6 ? dirty_109 : _GEN_6026; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7064 = _T_6 ? dirty_110 : _GEN_6027; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7065 = _T_6 ? dirty_111 : _GEN_6028; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7066 = _T_6 ? dirty_112 : _GEN_6029; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7067 = _T_6 ? dirty_113 : _GEN_6030; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7068 = _T_6 ? dirty_114 : _GEN_6031; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7069 = _T_6 ? dirty_115 : _GEN_6032; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7070 = _T_6 ? dirty_116 : _GEN_6033; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7071 = _T_6 ? dirty_117 : _GEN_6034; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7072 = _T_6 ? dirty_118 : _GEN_6035; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7073 = _T_6 ? dirty_119 : _GEN_6036; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7074 = _T_6 ? dirty_120 : _GEN_6037; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7075 = _T_6 ? dirty_121 : _GEN_6038; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7076 = _T_6 ? dirty_122 : _GEN_6039; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7077 = _T_6 ? dirty_123 : _GEN_6040; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7078 = _T_6 ? dirty_124 : _GEN_6041; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7079 = _T_6 ? dirty_125 : _GEN_6042; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7080 = _T_6 ? dirty_126 : _GEN_6043; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7081 = _T_6 ? dirty_127 : _GEN_6044; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7082 = _T_6 ? dirty_128 : _GEN_6045; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7083 = _T_6 ? dirty_129 : _GEN_6046; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7084 = _T_6 ? dirty_130 : _GEN_6047; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7085 = _T_6 ? dirty_131 : _GEN_6048; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7086 = _T_6 ? dirty_132 : _GEN_6049; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7087 = _T_6 ? dirty_133 : _GEN_6050; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7088 = _T_6 ? dirty_134 : _GEN_6051; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7089 = _T_6 ? dirty_135 : _GEN_6052; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7090 = _T_6 ? dirty_136 : _GEN_6053; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7091 = _T_6 ? dirty_137 : _GEN_6054; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7092 = _T_6 ? dirty_138 : _GEN_6055; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7093 = _T_6 ? dirty_139 : _GEN_6056; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7094 = _T_6 ? dirty_140 : _GEN_6057; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7095 = _T_6 ? dirty_141 : _GEN_6058; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7096 = _T_6 ? dirty_142 : _GEN_6059; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7097 = _T_6 ? dirty_143 : _GEN_6060; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7098 = _T_6 ? dirty_144 : _GEN_6061; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7099 = _T_6 ? dirty_145 : _GEN_6062; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7100 = _T_6 ? dirty_146 : _GEN_6063; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7101 = _T_6 ? dirty_147 : _GEN_6064; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7102 = _T_6 ? dirty_148 : _GEN_6065; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7103 = _T_6 ? dirty_149 : _GEN_6066; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7104 = _T_6 ? dirty_150 : _GEN_6067; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7105 = _T_6 ? dirty_151 : _GEN_6068; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7106 = _T_6 ? dirty_152 : _GEN_6069; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7107 = _T_6 ? dirty_153 : _GEN_6070; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7108 = _T_6 ? dirty_154 : _GEN_6071; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7109 = _T_6 ? dirty_155 : _GEN_6072; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7110 = _T_6 ? dirty_156 : _GEN_6073; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7111 = _T_6 ? dirty_157 : _GEN_6074; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7112 = _T_6 ? dirty_158 : _GEN_6075; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7113 = _T_6 ? dirty_159 : _GEN_6076; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7114 = _T_6 ? dirty_160 : _GEN_6077; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7115 = _T_6 ? dirty_161 : _GEN_6078; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7116 = _T_6 ? dirty_162 : _GEN_6079; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7117 = _T_6 ? dirty_163 : _GEN_6080; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7118 = _T_6 ? dirty_164 : _GEN_6081; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7119 = _T_6 ? dirty_165 : _GEN_6082; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7120 = _T_6 ? dirty_166 : _GEN_6083; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7121 = _T_6 ? dirty_167 : _GEN_6084; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7122 = _T_6 ? dirty_168 : _GEN_6085; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7123 = _T_6 ? dirty_169 : _GEN_6086; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7124 = _T_6 ? dirty_170 : _GEN_6087; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7125 = _T_6 ? dirty_171 : _GEN_6088; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7126 = _T_6 ? dirty_172 : _GEN_6089; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7127 = _T_6 ? dirty_173 : _GEN_6090; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7128 = _T_6 ? dirty_174 : _GEN_6091; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7129 = _T_6 ? dirty_175 : _GEN_6092; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7130 = _T_6 ? dirty_176 : _GEN_6093; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7131 = _T_6 ? dirty_177 : _GEN_6094; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7132 = _T_6 ? dirty_178 : _GEN_6095; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7133 = _T_6 ? dirty_179 : _GEN_6096; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7134 = _T_6 ? dirty_180 : _GEN_6097; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7135 = _T_6 ? dirty_181 : _GEN_6098; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7136 = _T_6 ? dirty_182 : _GEN_6099; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7137 = _T_6 ? dirty_183 : _GEN_6100; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7138 = _T_6 ? dirty_184 : _GEN_6101; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7139 = _T_6 ? dirty_185 : _GEN_6102; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7140 = _T_6 ? dirty_186 : _GEN_6103; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7141 = _T_6 ? dirty_187 : _GEN_6104; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7142 = _T_6 ? dirty_188 : _GEN_6105; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7143 = _T_6 ? dirty_189 : _GEN_6106; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7144 = _T_6 ? dirty_190 : _GEN_6107; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7145 = _T_6 ? dirty_191 : _GEN_6108; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7146 = _T_6 ? dirty_192 : _GEN_6109; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7147 = _T_6 ? dirty_193 : _GEN_6110; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7148 = _T_6 ? dirty_194 : _GEN_6111; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7149 = _T_6 ? dirty_195 : _GEN_6112; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7150 = _T_6 ? dirty_196 : _GEN_6113; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7151 = _T_6 ? dirty_197 : _GEN_6114; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7152 = _T_6 ? dirty_198 : _GEN_6115; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7153 = _T_6 ? dirty_199 : _GEN_6116; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7154 = _T_6 ? dirty_200 : _GEN_6117; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7155 = _T_6 ? dirty_201 : _GEN_6118; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7156 = _T_6 ? dirty_202 : _GEN_6119; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7157 = _T_6 ? dirty_203 : _GEN_6120; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7158 = _T_6 ? dirty_204 : _GEN_6121; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7159 = _T_6 ? dirty_205 : _GEN_6122; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7160 = _T_6 ? dirty_206 : _GEN_6123; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7161 = _T_6 ? dirty_207 : _GEN_6124; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7162 = _T_6 ? dirty_208 : _GEN_6125; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7163 = _T_6 ? dirty_209 : _GEN_6126; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7164 = _T_6 ? dirty_210 : _GEN_6127; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7165 = _T_6 ? dirty_211 : _GEN_6128; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7166 = _T_6 ? dirty_212 : _GEN_6129; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7167 = _T_6 ? dirty_213 : _GEN_6130; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7168 = _T_6 ? dirty_214 : _GEN_6131; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7169 = _T_6 ? dirty_215 : _GEN_6132; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7170 = _T_6 ? dirty_216 : _GEN_6133; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7171 = _T_6 ? dirty_217 : _GEN_6134; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7172 = _T_6 ? dirty_218 : _GEN_6135; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7173 = _T_6 ? dirty_219 : _GEN_6136; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7174 = _T_6 ? dirty_220 : _GEN_6137; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7175 = _T_6 ? dirty_221 : _GEN_6138; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7176 = _T_6 ? dirty_222 : _GEN_6139; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7177 = _T_6 ? dirty_223 : _GEN_6140; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7178 = _T_6 ? dirty_224 : _GEN_6141; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7179 = _T_6 ? dirty_225 : _GEN_6142; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7180 = _T_6 ? dirty_226 : _GEN_6143; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7181 = _T_6 ? dirty_227 : _GEN_6144; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7182 = _T_6 ? dirty_228 : _GEN_6145; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7183 = _T_6 ? dirty_229 : _GEN_6146; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7184 = _T_6 ? dirty_230 : _GEN_6147; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7185 = _T_6 ? dirty_231 : _GEN_6148; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7186 = _T_6 ? dirty_232 : _GEN_6149; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7187 = _T_6 ? dirty_233 : _GEN_6150; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7188 = _T_6 ? dirty_234 : _GEN_6151; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7189 = _T_6 ? dirty_235 : _GEN_6152; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7190 = _T_6 ? dirty_236 : _GEN_6153; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7191 = _T_6 ? dirty_237 : _GEN_6154; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7192 = _T_6 ? dirty_238 : _GEN_6155; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7193 = _T_6 ? dirty_239 : _GEN_6156; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7194 = _T_6 ? dirty_240 : _GEN_6157; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7195 = _T_6 ? dirty_241 : _GEN_6158; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7196 = _T_6 ? dirty_242 : _GEN_6159; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7197 = _T_6 ? dirty_243 : _GEN_6160; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7198 = _T_6 ? dirty_244 : _GEN_6161; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7199 = _T_6 ? dirty_245 : _GEN_6162; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7200 = _T_6 ? dirty_246 : _GEN_6163; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7201 = _T_6 ? dirty_247 : _GEN_6164; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7202 = _T_6 ? dirty_248 : _GEN_6165; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7203 = _T_6 ? dirty_249 : _GEN_6166; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7204 = _T_6 ? dirty_250 : _GEN_6167; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7205 = _T_6 ? dirty_251 : _GEN_6168; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7206 = _T_6 ? dirty_252 : _GEN_6169; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7207 = _T_6 ? dirty_253 : _GEN_6170; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7208 = _T_6 ? dirty_254 : _GEN_6171; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7209 = _T_6 ? dirty_255 : _GEN_6172; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire [3:0] _GEN_7210 = _T_6 ? offset_0 : _GEN_6173; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7211 = _T_6 ? offset_1 : _GEN_6174; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7212 = _T_6 ? offset_2 : _GEN_6175; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7213 = _T_6 ? offset_3 : _GEN_6176; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7214 = _T_6 ? offset_4 : _GEN_6177; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7215 = _T_6 ? offset_5 : _GEN_6178; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7216 = _T_6 ? offset_6 : _GEN_6179; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7217 = _T_6 ? offset_7 : _GEN_6180; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7218 = _T_6 ? offset_8 : _GEN_6181; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7219 = _T_6 ? offset_9 : _GEN_6182; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7220 = _T_6 ? offset_10 : _GEN_6183; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7221 = _T_6 ? offset_11 : _GEN_6184; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7222 = _T_6 ? offset_12 : _GEN_6185; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7223 = _T_6 ? offset_13 : _GEN_6186; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7224 = _T_6 ? offset_14 : _GEN_6187; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7225 = _T_6 ? offset_15 : _GEN_6188; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7226 = _T_6 ? offset_16 : _GEN_6189; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7227 = _T_6 ? offset_17 : _GEN_6190; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7228 = _T_6 ? offset_18 : _GEN_6191; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7229 = _T_6 ? offset_19 : _GEN_6192; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7230 = _T_6 ? offset_20 : _GEN_6193; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7231 = _T_6 ? offset_21 : _GEN_6194; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7232 = _T_6 ? offset_22 : _GEN_6195; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7233 = _T_6 ? offset_23 : _GEN_6196; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7234 = _T_6 ? offset_24 : _GEN_6197; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7235 = _T_6 ? offset_25 : _GEN_6198; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7236 = _T_6 ? offset_26 : _GEN_6199; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7237 = _T_6 ? offset_27 : _GEN_6200; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7238 = _T_6 ? offset_28 : _GEN_6201; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7239 = _T_6 ? offset_29 : _GEN_6202; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7240 = _T_6 ? offset_30 : _GEN_6203; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7241 = _T_6 ? offset_31 : _GEN_6204; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7242 = _T_6 ? offset_32 : _GEN_6205; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7243 = _T_6 ? offset_33 : _GEN_6206; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7244 = _T_6 ? offset_34 : _GEN_6207; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7245 = _T_6 ? offset_35 : _GEN_6208; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7246 = _T_6 ? offset_36 : _GEN_6209; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7247 = _T_6 ? offset_37 : _GEN_6210; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7248 = _T_6 ? offset_38 : _GEN_6211; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7249 = _T_6 ? offset_39 : _GEN_6212; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7250 = _T_6 ? offset_40 : _GEN_6213; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7251 = _T_6 ? offset_41 : _GEN_6214; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7252 = _T_6 ? offset_42 : _GEN_6215; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7253 = _T_6 ? offset_43 : _GEN_6216; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7254 = _T_6 ? offset_44 : _GEN_6217; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7255 = _T_6 ? offset_45 : _GEN_6218; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7256 = _T_6 ? offset_46 : _GEN_6219; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7257 = _T_6 ? offset_47 : _GEN_6220; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7258 = _T_6 ? offset_48 : _GEN_6221; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7259 = _T_6 ? offset_49 : _GEN_6222; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7260 = _T_6 ? offset_50 : _GEN_6223; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7261 = _T_6 ? offset_51 : _GEN_6224; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7262 = _T_6 ? offset_52 : _GEN_6225; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7263 = _T_6 ? offset_53 : _GEN_6226; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7264 = _T_6 ? offset_54 : _GEN_6227; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7265 = _T_6 ? offset_55 : _GEN_6228; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7266 = _T_6 ? offset_56 : _GEN_6229; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7267 = _T_6 ? offset_57 : _GEN_6230; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7268 = _T_6 ? offset_58 : _GEN_6231; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7269 = _T_6 ? offset_59 : _GEN_6232; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7270 = _T_6 ? offset_60 : _GEN_6233; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7271 = _T_6 ? offset_61 : _GEN_6234; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7272 = _T_6 ? offset_62 : _GEN_6235; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7273 = _T_6 ? offset_63 : _GEN_6236; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7274 = _T_6 ? offset_64 : _GEN_6237; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7275 = _T_6 ? offset_65 : _GEN_6238; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7276 = _T_6 ? offset_66 : _GEN_6239; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7277 = _T_6 ? offset_67 : _GEN_6240; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7278 = _T_6 ? offset_68 : _GEN_6241; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7279 = _T_6 ? offset_69 : _GEN_6242; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7280 = _T_6 ? offset_70 : _GEN_6243; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7281 = _T_6 ? offset_71 : _GEN_6244; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7282 = _T_6 ? offset_72 : _GEN_6245; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7283 = _T_6 ? offset_73 : _GEN_6246; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7284 = _T_6 ? offset_74 : _GEN_6247; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7285 = _T_6 ? offset_75 : _GEN_6248; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7286 = _T_6 ? offset_76 : _GEN_6249; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7287 = _T_6 ? offset_77 : _GEN_6250; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7288 = _T_6 ? offset_78 : _GEN_6251; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7289 = _T_6 ? offset_79 : _GEN_6252; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7290 = _T_6 ? offset_80 : _GEN_6253; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7291 = _T_6 ? offset_81 : _GEN_6254; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7292 = _T_6 ? offset_82 : _GEN_6255; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7293 = _T_6 ? offset_83 : _GEN_6256; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7294 = _T_6 ? offset_84 : _GEN_6257; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7295 = _T_6 ? offset_85 : _GEN_6258; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7296 = _T_6 ? offset_86 : _GEN_6259; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7297 = _T_6 ? offset_87 : _GEN_6260; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7298 = _T_6 ? offset_88 : _GEN_6261; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7299 = _T_6 ? offset_89 : _GEN_6262; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7300 = _T_6 ? offset_90 : _GEN_6263; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7301 = _T_6 ? offset_91 : _GEN_6264; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7302 = _T_6 ? offset_92 : _GEN_6265; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7303 = _T_6 ? offset_93 : _GEN_6266; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7304 = _T_6 ? offset_94 : _GEN_6267; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7305 = _T_6 ? offset_95 : _GEN_6268; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7306 = _T_6 ? offset_96 : _GEN_6269; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7307 = _T_6 ? offset_97 : _GEN_6270; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7308 = _T_6 ? offset_98 : _GEN_6271; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7309 = _T_6 ? offset_99 : _GEN_6272; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7310 = _T_6 ? offset_100 : _GEN_6273; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7311 = _T_6 ? offset_101 : _GEN_6274; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7312 = _T_6 ? offset_102 : _GEN_6275; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7313 = _T_6 ? offset_103 : _GEN_6276; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7314 = _T_6 ? offset_104 : _GEN_6277; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7315 = _T_6 ? offset_105 : _GEN_6278; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7316 = _T_6 ? offset_106 : _GEN_6279; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7317 = _T_6 ? offset_107 : _GEN_6280; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7318 = _T_6 ? offset_108 : _GEN_6281; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7319 = _T_6 ? offset_109 : _GEN_6282; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7320 = _T_6 ? offset_110 : _GEN_6283; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7321 = _T_6 ? offset_111 : _GEN_6284; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7322 = _T_6 ? offset_112 : _GEN_6285; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7323 = _T_6 ? offset_113 : _GEN_6286; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7324 = _T_6 ? offset_114 : _GEN_6287; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7325 = _T_6 ? offset_115 : _GEN_6288; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7326 = _T_6 ? offset_116 : _GEN_6289; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7327 = _T_6 ? offset_117 : _GEN_6290; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7328 = _T_6 ? offset_118 : _GEN_6291; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7329 = _T_6 ? offset_119 : _GEN_6292; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7330 = _T_6 ? offset_120 : _GEN_6293; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7331 = _T_6 ? offset_121 : _GEN_6294; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7332 = _T_6 ? offset_122 : _GEN_6295; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7333 = _T_6 ? offset_123 : _GEN_6296; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7334 = _T_6 ? offset_124 : _GEN_6297; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7335 = _T_6 ? offset_125 : _GEN_6298; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7336 = _T_6 ? offset_126 : _GEN_6299; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7337 = _T_6 ? offset_127 : _GEN_6300; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7338 = _T_6 ? offset_128 : _GEN_6301; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7339 = _T_6 ? offset_129 : _GEN_6302; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7340 = _T_6 ? offset_130 : _GEN_6303; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7341 = _T_6 ? offset_131 : _GEN_6304; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7342 = _T_6 ? offset_132 : _GEN_6305; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7343 = _T_6 ? offset_133 : _GEN_6306; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7344 = _T_6 ? offset_134 : _GEN_6307; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7345 = _T_6 ? offset_135 : _GEN_6308; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7346 = _T_6 ? offset_136 : _GEN_6309; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7347 = _T_6 ? offset_137 : _GEN_6310; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7348 = _T_6 ? offset_138 : _GEN_6311; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7349 = _T_6 ? offset_139 : _GEN_6312; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7350 = _T_6 ? offset_140 : _GEN_6313; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7351 = _T_6 ? offset_141 : _GEN_6314; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7352 = _T_6 ? offset_142 : _GEN_6315; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7353 = _T_6 ? offset_143 : _GEN_6316; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7354 = _T_6 ? offset_144 : _GEN_6317; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7355 = _T_6 ? offset_145 : _GEN_6318; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7356 = _T_6 ? offset_146 : _GEN_6319; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7357 = _T_6 ? offset_147 : _GEN_6320; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7358 = _T_6 ? offset_148 : _GEN_6321; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7359 = _T_6 ? offset_149 : _GEN_6322; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7360 = _T_6 ? offset_150 : _GEN_6323; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7361 = _T_6 ? offset_151 : _GEN_6324; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7362 = _T_6 ? offset_152 : _GEN_6325; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7363 = _T_6 ? offset_153 : _GEN_6326; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7364 = _T_6 ? offset_154 : _GEN_6327; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7365 = _T_6 ? offset_155 : _GEN_6328; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7366 = _T_6 ? offset_156 : _GEN_6329; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7367 = _T_6 ? offset_157 : _GEN_6330; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7368 = _T_6 ? offset_158 : _GEN_6331; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7369 = _T_6 ? offset_159 : _GEN_6332; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7370 = _T_6 ? offset_160 : _GEN_6333; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7371 = _T_6 ? offset_161 : _GEN_6334; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7372 = _T_6 ? offset_162 : _GEN_6335; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7373 = _T_6 ? offset_163 : _GEN_6336; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7374 = _T_6 ? offset_164 : _GEN_6337; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7375 = _T_6 ? offset_165 : _GEN_6338; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7376 = _T_6 ? offset_166 : _GEN_6339; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7377 = _T_6 ? offset_167 : _GEN_6340; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7378 = _T_6 ? offset_168 : _GEN_6341; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7379 = _T_6 ? offset_169 : _GEN_6342; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7380 = _T_6 ? offset_170 : _GEN_6343; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7381 = _T_6 ? offset_171 : _GEN_6344; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7382 = _T_6 ? offset_172 : _GEN_6345; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7383 = _T_6 ? offset_173 : _GEN_6346; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7384 = _T_6 ? offset_174 : _GEN_6347; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7385 = _T_6 ? offset_175 : _GEN_6348; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7386 = _T_6 ? offset_176 : _GEN_6349; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7387 = _T_6 ? offset_177 : _GEN_6350; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7388 = _T_6 ? offset_178 : _GEN_6351; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7389 = _T_6 ? offset_179 : _GEN_6352; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7390 = _T_6 ? offset_180 : _GEN_6353; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7391 = _T_6 ? offset_181 : _GEN_6354; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7392 = _T_6 ? offset_182 : _GEN_6355; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7393 = _T_6 ? offset_183 : _GEN_6356; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7394 = _T_6 ? offset_184 : _GEN_6357; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7395 = _T_6 ? offset_185 : _GEN_6358; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7396 = _T_6 ? offset_186 : _GEN_6359; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7397 = _T_6 ? offset_187 : _GEN_6360; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7398 = _T_6 ? offset_188 : _GEN_6361; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7399 = _T_6 ? offset_189 : _GEN_6362; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7400 = _T_6 ? offset_190 : _GEN_6363; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7401 = _T_6 ? offset_191 : _GEN_6364; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7402 = _T_6 ? offset_192 : _GEN_6365; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7403 = _T_6 ? offset_193 : _GEN_6366; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7404 = _T_6 ? offset_194 : _GEN_6367; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7405 = _T_6 ? offset_195 : _GEN_6368; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7406 = _T_6 ? offset_196 : _GEN_6369; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7407 = _T_6 ? offset_197 : _GEN_6370; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7408 = _T_6 ? offset_198 : _GEN_6371; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7409 = _T_6 ? offset_199 : _GEN_6372; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7410 = _T_6 ? offset_200 : _GEN_6373; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7411 = _T_6 ? offset_201 : _GEN_6374; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7412 = _T_6 ? offset_202 : _GEN_6375; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7413 = _T_6 ? offset_203 : _GEN_6376; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7414 = _T_6 ? offset_204 : _GEN_6377; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7415 = _T_6 ? offset_205 : _GEN_6378; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7416 = _T_6 ? offset_206 : _GEN_6379; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7417 = _T_6 ? offset_207 : _GEN_6380; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7418 = _T_6 ? offset_208 : _GEN_6381; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7419 = _T_6 ? offset_209 : _GEN_6382; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7420 = _T_6 ? offset_210 : _GEN_6383; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7421 = _T_6 ? offset_211 : _GEN_6384; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7422 = _T_6 ? offset_212 : _GEN_6385; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7423 = _T_6 ? offset_213 : _GEN_6386; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7424 = _T_6 ? offset_214 : _GEN_6387; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7425 = _T_6 ? offset_215 : _GEN_6388; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7426 = _T_6 ? offset_216 : _GEN_6389; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7427 = _T_6 ? offset_217 : _GEN_6390; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7428 = _T_6 ? offset_218 : _GEN_6391; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7429 = _T_6 ? offset_219 : _GEN_6392; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7430 = _T_6 ? offset_220 : _GEN_6393; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7431 = _T_6 ? offset_221 : _GEN_6394; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7432 = _T_6 ? offset_222 : _GEN_6395; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7433 = _T_6 ? offset_223 : _GEN_6396; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7434 = _T_6 ? offset_224 : _GEN_6397; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7435 = _T_6 ? offset_225 : _GEN_6398; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7436 = _T_6 ? offset_226 : _GEN_6399; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7437 = _T_6 ? offset_227 : _GEN_6400; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7438 = _T_6 ? offset_228 : _GEN_6401; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7439 = _T_6 ? offset_229 : _GEN_6402; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7440 = _T_6 ? offset_230 : _GEN_6403; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7441 = _T_6 ? offset_231 : _GEN_6404; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7442 = _T_6 ? offset_232 : _GEN_6405; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7443 = _T_6 ? offset_233 : _GEN_6406; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7444 = _T_6 ? offset_234 : _GEN_6407; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7445 = _T_6 ? offset_235 : _GEN_6408; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7446 = _T_6 ? offset_236 : _GEN_6409; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7447 = _T_6 ? offset_237 : _GEN_6410; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7448 = _T_6 ? offset_238 : _GEN_6411; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7449 = _T_6 ? offset_239 : _GEN_6412; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7450 = _T_6 ? offset_240 : _GEN_6413; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7451 = _T_6 ? offset_241 : _GEN_6414; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7452 = _T_6 ? offset_242 : _GEN_6415; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7453 = _T_6 ? offset_243 : _GEN_6416; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7454 = _T_6 ? offset_244 : _GEN_6417; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7455 = _T_6 ? offset_245 : _GEN_6418; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7456 = _T_6 ? offset_246 : _GEN_6419; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7457 = _T_6 ? offset_247 : _GEN_6420; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7458 = _T_6 ? offset_248 : _GEN_6421; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7459 = _T_6 ? offset_249 : _GEN_6422; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7460 = _T_6 ? offset_250 : _GEN_6423; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7461 = _T_6 ? offset_251 : _GEN_6424; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7462 = _T_6 ? offset_252 : _GEN_6425; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7463 = _T_6 ? offset_253 : _GEN_6426; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7464 = _T_6 ? offset_254 : _GEN_6427; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7465 = _T_6 ? offset_255 : _GEN_6428; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [2:0] _GEN_7466 = _T_5 ? 3'h4 : _GEN_6430; // @[Conditional.scala 39:67 Dcache.scala 173:15]
  wire [31:0] _GEN_7467 = _T_5 ? 32'h0 : _GEN_6431; // @[Conditional.scala 39:67]
  wire  _GEN_7471 = _T_5 ? 1'h0 : _T_6 & _GEN_4377; // @[Conditional.scala 39:67]
  wire  _GEN_7473 = _T_5 ? cache_fill : _GEN_6437; // @[Conditional.scala 39:67 Dcache.scala 116:28]
  wire  _GEN_7474 = _T_5 ? cache_wen : _GEN_6438; // @[Conditional.scala 39:67 Dcache.scala 117:28]
  wire [127:0] _GEN_7475 = _T_5 ? cache_wdata : _GEN_6439; // @[Conditional.scala 39:67 Dcache.scala 118:28]
  wire [127:0] _GEN_7476 = _T_5 ? cache_strb : _GEN_6440; // @[Conditional.scala 39:67 Dcache.scala 119:28]
  wire  _GEN_7477 = _T_5 ? data_ready : _GEN_6441; // @[Conditional.scala 39:67 Dcache.scala 46:28]
  wire  _GEN_7478 = _T_5 ? valid_0 : _GEN_6442; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7479 = _T_5 ? valid_1 : _GEN_6443; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7480 = _T_5 ? valid_2 : _GEN_6444; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7481 = _T_5 ? valid_3 : _GEN_6445; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7482 = _T_5 ? valid_4 : _GEN_6446; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7483 = _T_5 ? valid_5 : _GEN_6447; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7484 = _T_5 ? valid_6 : _GEN_6448; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7485 = _T_5 ? valid_7 : _GEN_6449; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7486 = _T_5 ? valid_8 : _GEN_6450; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7487 = _T_5 ? valid_9 : _GEN_6451; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7488 = _T_5 ? valid_10 : _GEN_6452; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7489 = _T_5 ? valid_11 : _GEN_6453; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7490 = _T_5 ? valid_12 : _GEN_6454; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7491 = _T_5 ? valid_13 : _GEN_6455; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7492 = _T_5 ? valid_14 : _GEN_6456; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7493 = _T_5 ? valid_15 : _GEN_6457; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7494 = _T_5 ? valid_16 : _GEN_6458; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7495 = _T_5 ? valid_17 : _GEN_6459; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7496 = _T_5 ? valid_18 : _GEN_6460; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7497 = _T_5 ? valid_19 : _GEN_6461; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7498 = _T_5 ? valid_20 : _GEN_6462; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7499 = _T_5 ? valid_21 : _GEN_6463; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7500 = _T_5 ? valid_22 : _GEN_6464; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7501 = _T_5 ? valid_23 : _GEN_6465; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7502 = _T_5 ? valid_24 : _GEN_6466; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7503 = _T_5 ? valid_25 : _GEN_6467; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7504 = _T_5 ? valid_26 : _GEN_6468; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7505 = _T_5 ? valid_27 : _GEN_6469; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7506 = _T_5 ? valid_28 : _GEN_6470; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7507 = _T_5 ? valid_29 : _GEN_6471; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7508 = _T_5 ? valid_30 : _GEN_6472; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7509 = _T_5 ? valid_31 : _GEN_6473; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7510 = _T_5 ? valid_32 : _GEN_6474; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7511 = _T_5 ? valid_33 : _GEN_6475; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7512 = _T_5 ? valid_34 : _GEN_6476; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7513 = _T_5 ? valid_35 : _GEN_6477; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7514 = _T_5 ? valid_36 : _GEN_6478; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7515 = _T_5 ? valid_37 : _GEN_6479; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7516 = _T_5 ? valid_38 : _GEN_6480; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7517 = _T_5 ? valid_39 : _GEN_6481; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7518 = _T_5 ? valid_40 : _GEN_6482; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7519 = _T_5 ? valid_41 : _GEN_6483; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7520 = _T_5 ? valid_42 : _GEN_6484; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7521 = _T_5 ? valid_43 : _GEN_6485; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7522 = _T_5 ? valid_44 : _GEN_6486; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7523 = _T_5 ? valid_45 : _GEN_6487; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7524 = _T_5 ? valid_46 : _GEN_6488; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7525 = _T_5 ? valid_47 : _GEN_6489; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7526 = _T_5 ? valid_48 : _GEN_6490; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7527 = _T_5 ? valid_49 : _GEN_6491; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7528 = _T_5 ? valid_50 : _GEN_6492; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7529 = _T_5 ? valid_51 : _GEN_6493; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7530 = _T_5 ? valid_52 : _GEN_6494; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7531 = _T_5 ? valid_53 : _GEN_6495; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7532 = _T_5 ? valid_54 : _GEN_6496; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7533 = _T_5 ? valid_55 : _GEN_6497; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7534 = _T_5 ? valid_56 : _GEN_6498; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7535 = _T_5 ? valid_57 : _GEN_6499; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7536 = _T_5 ? valid_58 : _GEN_6500; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7537 = _T_5 ? valid_59 : _GEN_6501; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7538 = _T_5 ? valid_60 : _GEN_6502; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7539 = _T_5 ? valid_61 : _GEN_6503; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7540 = _T_5 ? valid_62 : _GEN_6504; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7541 = _T_5 ? valid_63 : _GEN_6505; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7542 = _T_5 ? valid_64 : _GEN_6506; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7543 = _T_5 ? valid_65 : _GEN_6507; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7544 = _T_5 ? valid_66 : _GEN_6508; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7545 = _T_5 ? valid_67 : _GEN_6509; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7546 = _T_5 ? valid_68 : _GEN_6510; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7547 = _T_5 ? valid_69 : _GEN_6511; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7548 = _T_5 ? valid_70 : _GEN_6512; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7549 = _T_5 ? valid_71 : _GEN_6513; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7550 = _T_5 ? valid_72 : _GEN_6514; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7551 = _T_5 ? valid_73 : _GEN_6515; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7552 = _T_5 ? valid_74 : _GEN_6516; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7553 = _T_5 ? valid_75 : _GEN_6517; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7554 = _T_5 ? valid_76 : _GEN_6518; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7555 = _T_5 ? valid_77 : _GEN_6519; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7556 = _T_5 ? valid_78 : _GEN_6520; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7557 = _T_5 ? valid_79 : _GEN_6521; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7558 = _T_5 ? valid_80 : _GEN_6522; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7559 = _T_5 ? valid_81 : _GEN_6523; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7560 = _T_5 ? valid_82 : _GEN_6524; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7561 = _T_5 ? valid_83 : _GEN_6525; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7562 = _T_5 ? valid_84 : _GEN_6526; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7563 = _T_5 ? valid_85 : _GEN_6527; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7564 = _T_5 ? valid_86 : _GEN_6528; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7565 = _T_5 ? valid_87 : _GEN_6529; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7566 = _T_5 ? valid_88 : _GEN_6530; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7567 = _T_5 ? valid_89 : _GEN_6531; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7568 = _T_5 ? valid_90 : _GEN_6532; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7569 = _T_5 ? valid_91 : _GEN_6533; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7570 = _T_5 ? valid_92 : _GEN_6534; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7571 = _T_5 ? valid_93 : _GEN_6535; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7572 = _T_5 ? valid_94 : _GEN_6536; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7573 = _T_5 ? valid_95 : _GEN_6537; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7574 = _T_5 ? valid_96 : _GEN_6538; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7575 = _T_5 ? valid_97 : _GEN_6539; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7576 = _T_5 ? valid_98 : _GEN_6540; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7577 = _T_5 ? valid_99 : _GEN_6541; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7578 = _T_5 ? valid_100 : _GEN_6542; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7579 = _T_5 ? valid_101 : _GEN_6543; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7580 = _T_5 ? valid_102 : _GEN_6544; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7581 = _T_5 ? valid_103 : _GEN_6545; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7582 = _T_5 ? valid_104 : _GEN_6546; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7583 = _T_5 ? valid_105 : _GEN_6547; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7584 = _T_5 ? valid_106 : _GEN_6548; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7585 = _T_5 ? valid_107 : _GEN_6549; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7586 = _T_5 ? valid_108 : _GEN_6550; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7587 = _T_5 ? valid_109 : _GEN_6551; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7588 = _T_5 ? valid_110 : _GEN_6552; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7589 = _T_5 ? valid_111 : _GEN_6553; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7590 = _T_5 ? valid_112 : _GEN_6554; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7591 = _T_5 ? valid_113 : _GEN_6555; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7592 = _T_5 ? valid_114 : _GEN_6556; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7593 = _T_5 ? valid_115 : _GEN_6557; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7594 = _T_5 ? valid_116 : _GEN_6558; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7595 = _T_5 ? valid_117 : _GEN_6559; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7596 = _T_5 ? valid_118 : _GEN_6560; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7597 = _T_5 ? valid_119 : _GEN_6561; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7598 = _T_5 ? valid_120 : _GEN_6562; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7599 = _T_5 ? valid_121 : _GEN_6563; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7600 = _T_5 ? valid_122 : _GEN_6564; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7601 = _T_5 ? valid_123 : _GEN_6565; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7602 = _T_5 ? valid_124 : _GEN_6566; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7603 = _T_5 ? valid_125 : _GEN_6567; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7604 = _T_5 ? valid_126 : _GEN_6568; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7605 = _T_5 ? valid_127 : _GEN_6569; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7606 = _T_5 ? valid_128 : _GEN_6570; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7607 = _T_5 ? valid_129 : _GEN_6571; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7608 = _T_5 ? valid_130 : _GEN_6572; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7609 = _T_5 ? valid_131 : _GEN_6573; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7610 = _T_5 ? valid_132 : _GEN_6574; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7611 = _T_5 ? valid_133 : _GEN_6575; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7612 = _T_5 ? valid_134 : _GEN_6576; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7613 = _T_5 ? valid_135 : _GEN_6577; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7614 = _T_5 ? valid_136 : _GEN_6578; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7615 = _T_5 ? valid_137 : _GEN_6579; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7616 = _T_5 ? valid_138 : _GEN_6580; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7617 = _T_5 ? valid_139 : _GEN_6581; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7618 = _T_5 ? valid_140 : _GEN_6582; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7619 = _T_5 ? valid_141 : _GEN_6583; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7620 = _T_5 ? valid_142 : _GEN_6584; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7621 = _T_5 ? valid_143 : _GEN_6585; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7622 = _T_5 ? valid_144 : _GEN_6586; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7623 = _T_5 ? valid_145 : _GEN_6587; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7624 = _T_5 ? valid_146 : _GEN_6588; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7625 = _T_5 ? valid_147 : _GEN_6589; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7626 = _T_5 ? valid_148 : _GEN_6590; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7627 = _T_5 ? valid_149 : _GEN_6591; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7628 = _T_5 ? valid_150 : _GEN_6592; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7629 = _T_5 ? valid_151 : _GEN_6593; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7630 = _T_5 ? valid_152 : _GEN_6594; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7631 = _T_5 ? valid_153 : _GEN_6595; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7632 = _T_5 ? valid_154 : _GEN_6596; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7633 = _T_5 ? valid_155 : _GEN_6597; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7634 = _T_5 ? valid_156 : _GEN_6598; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7635 = _T_5 ? valid_157 : _GEN_6599; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7636 = _T_5 ? valid_158 : _GEN_6600; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7637 = _T_5 ? valid_159 : _GEN_6601; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7638 = _T_5 ? valid_160 : _GEN_6602; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7639 = _T_5 ? valid_161 : _GEN_6603; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7640 = _T_5 ? valid_162 : _GEN_6604; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7641 = _T_5 ? valid_163 : _GEN_6605; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7642 = _T_5 ? valid_164 : _GEN_6606; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7643 = _T_5 ? valid_165 : _GEN_6607; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7644 = _T_5 ? valid_166 : _GEN_6608; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7645 = _T_5 ? valid_167 : _GEN_6609; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7646 = _T_5 ? valid_168 : _GEN_6610; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7647 = _T_5 ? valid_169 : _GEN_6611; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7648 = _T_5 ? valid_170 : _GEN_6612; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7649 = _T_5 ? valid_171 : _GEN_6613; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7650 = _T_5 ? valid_172 : _GEN_6614; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7651 = _T_5 ? valid_173 : _GEN_6615; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7652 = _T_5 ? valid_174 : _GEN_6616; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7653 = _T_5 ? valid_175 : _GEN_6617; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7654 = _T_5 ? valid_176 : _GEN_6618; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7655 = _T_5 ? valid_177 : _GEN_6619; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7656 = _T_5 ? valid_178 : _GEN_6620; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7657 = _T_5 ? valid_179 : _GEN_6621; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7658 = _T_5 ? valid_180 : _GEN_6622; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7659 = _T_5 ? valid_181 : _GEN_6623; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7660 = _T_5 ? valid_182 : _GEN_6624; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7661 = _T_5 ? valid_183 : _GEN_6625; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7662 = _T_5 ? valid_184 : _GEN_6626; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7663 = _T_5 ? valid_185 : _GEN_6627; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7664 = _T_5 ? valid_186 : _GEN_6628; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7665 = _T_5 ? valid_187 : _GEN_6629; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7666 = _T_5 ? valid_188 : _GEN_6630; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7667 = _T_5 ? valid_189 : _GEN_6631; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7668 = _T_5 ? valid_190 : _GEN_6632; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7669 = _T_5 ? valid_191 : _GEN_6633; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7670 = _T_5 ? valid_192 : _GEN_6634; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7671 = _T_5 ? valid_193 : _GEN_6635; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7672 = _T_5 ? valid_194 : _GEN_6636; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7673 = _T_5 ? valid_195 : _GEN_6637; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7674 = _T_5 ? valid_196 : _GEN_6638; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7675 = _T_5 ? valid_197 : _GEN_6639; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7676 = _T_5 ? valid_198 : _GEN_6640; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7677 = _T_5 ? valid_199 : _GEN_6641; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7678 = _T_5 ? valid_200 : _GEN_6642; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7679 = _T_5 ? valid_201 : _GEN_6643; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7680 = _T_5 ? valid_202 : _GEN_6644; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7681 = _T_5 ? valid_203 : _GEN_6645; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7682 = _T_5 ? valid_204 : _GEN_6646; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7683 = _T_5 ? valid_205 : _GEN_6647; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7684 = _T_5 ? valid_206 : _GEN_6648; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7685 = _T_5 ? valid_207 : _GEN_6649; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7686 = _T_5 ? valid_208 : _GEN_6650; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7687 = _T_5 ? valid_209 : _GEN_6651; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7688 = _T_5 ? valid_210 : _GEN_6652; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7689 = _T_5 ? valid_211 : _GEN_6653; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7690 = _T_5 ? valid_212 : _GEN_6654; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7691 = _T_5 ? valid_213 : _GEN_6655; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7692 = _T_5 ? valid_214 : _GEN_6656; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7693 = _T_5 ? valid_215 : _GEN_6657; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7694 = _T_5 ? valid_216 : _GEN_6658; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7695 = _T_5 ? valid_217 : _GEN_6659; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7696 = _T_5 ? valid_218 : _GEN_6660; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7697 = _T_5 ? valid_219 : _GEN_6661; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7698 = _T_5 ? valid_220 : _GEN_6662; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7699 = _T_5 ? valid_221 : _GEN_6663; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7700 = _T_5 ? valid_222 : _GEN_6664; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7701 = _T_5 ? valid_223 : _GEN_6665; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7702 = _T_5 ? valid_224 : _GEN_6666; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7703 = _T_5 ? valid_225 : _GEN_6667; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7704 = _T_5 ? valid_226 : _GEN_6668; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7705 = _T_5 ? valid_227 : _GEN_6669; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7706 = _T_5 ? valid_228 : _GEN_6670; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7707 = _T_5 ? valid_229 : _GEN_6671; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7708 = _T_5 ? valid_230 : _GEN_6672; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7709 = _T_5 ? valid_231 : _GEN_6673; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7710 = _T_5 ? valid_232 : _GEN_6674; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7711 = _T_5 ? valid_233 : _GEN_6675; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7712 = _T_5 ? valid_234 : _GEN_6676; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7713 = _T_5 ? valid_235 : _GEN_6677; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7714 = _T_5 ? valid_236 : _GEN_6678; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7715 = _T_5 ? valid_237 : _GEN_6679; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7716 = _T_5 ? valid_238 : _GEN_6680; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7717 = _T_5 ? valid_239 : _GEN_6681; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7718 = _T_5 ? valid_240 : _GEN_6682; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7719 = _T_5 ? valid_241 : _GEN_6683; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7720 = _T_5 ? valid_242 : _GEN_6684; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7721 = _T_5 ? valid_243 : _GEN_6685; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7722 = _T_5 ? valid_244 : _GEN_6686; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7723 = _T_5 ? valid_245 : _GEN_6687; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7724 = _T_5 ? valid_246 : _GEN_6688; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7725 = _T_5 ? valid_247 : _GEN_6689; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7726 = _T_5 ? valid_248 : _GEN_6690; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7727 = _T_5 ? valid_249 : _GEN_6691; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7728 = _T_5 ? valid_250 : _GEN_6692; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7729 = _T_5 ? valid_251 : _GEN_6693; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7730 = _T_5 ? valid_252 : _GEN_6694; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7731 = _T_5 ? valid_253 : _GEN_6695; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7732 = _T_5 ? valid_254 : _GEN_6696; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_7733 = _T_5 ? valid_255 : _GEN_6697; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire [19:0] _GEN_7734 = _T_5 ? tag_0 : _GEN_6698; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7735 = _T_5 ? tag_1 : _GEN_6699; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7736 = _T_5 ? tag_2 : _GEN_6700; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7737 = _T_5 ? tag_3 : _GEN_6701; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7738 = _T_5 ? tag_4 : _GEN_6702; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7739 = _T_5 ? tag_5 : _GEN_6703; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7740 = _T_5 ? tag_6 : _GEN_6704; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7741 = _T_5 ? tag_7 : _GEN_6705; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7742 = _T_5 ? tag_8 : _GEN_6706; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7743 = _T_5 ? tag_9 : _GEN_6707; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7744 = _T_5 ? tag_10 : _GEN_6708; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7745 = _T_5 ? tag_11 : _GEN_6709; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7746 = _T_5 ? tag_12 : _GEN_6710; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7747 = _T_5 ? tag_13 : _GEN_6711; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7748 = _T_5 ? tag_14 : _GEN_6712; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7749 = _T_5 ? tag_15 : _GEN_6713; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7750 = _T_5 ? tag_16 : _GEN_6714; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7751 = _T_5 ? tag_17 : _GEN_6715; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7752 = _T_5 ? tag_18 : _GEN_6716; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7753 = _T_5 ? tag_19 : _GEN_6717; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7754 = _T_5 ? tag_20 : _GEN_6718; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7755 = _T_5 ? tag_21 : _GEN_6719; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7756 = _T_5 ? tag_22 : _GEN_6720; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7757 = _T_5 ? tag_23 : _GEN_6721; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7758 = _T_5 ? tag_24 : _GEN_6722; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7759 = _T_5 ? tag_25 : _GEN_6723; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7760 = _T_5 ? tag_26 : _GEN_6724; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7761 = _T_5 ? tag_27 : _GEN_6725; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7762 = _T_5 ? tag_28 : _GEN_6726; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7763 = _T_5 ? tag_29 : _GEN_6727; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7764 = _T_5 ? tag_30 : _GEN_6728; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7765 = _T_5 ? tag_31 : _GEN_6729; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7766 = _T_5 ? tag_32 : _GEN_6730; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7767 = _T_5 ? tag_33 : _GEN_6731; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7768 = _T_5 ? tag_34 : _GEN_6732; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7769 = _T_5 ? tag_35 : _GEN_6733; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7770 = _T_5 ? tag_36 : _GEN_6734; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7771 = _T_5 ? tag_37 : _GEN_6735; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7772 = _T_5 ? tag_38 : _GEN_6736; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7773 = _T_5 ? tag_39 : _GEN_6737; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7774 = _T_5 ? tag_40 : _GEN_6738; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7775 = _T_5 ? tag_41 : _GEN_6739; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7776 = _T_5 ? tag_42 : _GEN_6740; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7777 = _T_5 ? tag_43 : _GEN_6741; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7778 = _T_5 ? tag_44 : _GEN_6742; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7779 = _T_5 ? tag_45 : _GEN_6743; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7780 = _T_5 ? tag_46 : _GEN_6744; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7781 = _T_5 ? tag_47 : _GEN_6745; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7782 = _T_5 ? tag_48 : _GEN_6746; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7783 = _T_5 ? tag_49 : _GEN_6747; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7784 = _T_5 ? tag_50 : _GEN_6748; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7785 = _T_5 ? tag_51 : _GEN_6749; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7786 = _T_5 ? tag_52 : _GEN_6750; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7787 = _T_5 ? tag_53 : _GEN_6751; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7788 = _T_5 ? tag_54 : _GEN_6752; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7789 = _T_5 ? tag_55 : _GEN_6753; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7790 = _T_5 ? tag_56 : _GEN_6754; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7791 = _T_5 ? tag_57 : _GEN_6755; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7792 = _T_5 ? tag_58 : _GEN_6756; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7793 = _T_5 ? tag_59 : _GEN_6757; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7794 = _T_5 ? tag_60 : _GEN_6758; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7795 = _T_5 ? tag_61 : _GEN_6759; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7796 = _T_5 ? tag_62 : _GEN_6760; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7797 = _T_5 ? tag_63 : _GEN_6761; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7798 = _T_5 ? tag_64 : _GEN_6762; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7799 = _T_5 ? tag_65 : _GEN_6763; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7800 = _T_5 ? tag_66 : _GEN_6764; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7801 = _T_5 ? tag_67 : _GEN_6765; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7802 = _T_5 ? tag_68 : _GEN_6766; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7803 = _T_5 ? tag_69 : _GEN_6767; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7804 = _T_5 ? tag_70 : _GEN_6768; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7805 = _T_5 ? tag_71 : _GEN_6769; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7806 = _T_5 ? tag_72 : _GEN_6770; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7807 = _T_5 ? tag_73 : _GEN_6771; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7808 = _T_5 ? tag_74 : _GEN_6772; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7809 = _T_5 ? tag_75 : _GEN_6773; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7810 = _T_5 ? tag_76 : _GEN_6774; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7811 = _T_5 ? tag_77 : _GEN_6775; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7812 = _T_5 ? tag_78 : _GEN_6776; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7813 = _T_5 ? tag_79 : _GEN_6777; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7814 = _T_5 ? tag_80 : _GEN_6778; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7815 = _T_5 ? tag_81 : _GEN_6779; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7816 = _T_5 ? tag_82 : _GEN_6780; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7817 = _T_5 ? tag_83 : _GEN_6781; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7818 = _T_5 ? tag_84 : _GEN_6782; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7819 = _T_5 ? tag_85 : _GEN_6783; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7820 = _T_5 ? tag_86 : _GEN_6784; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7821 = _T_5 ? tag_87 : _GEN_6785; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7822 = _T_5 ? tag_88 : _GEN_6786; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7823 = _T_5 ? tag_89 : _GEN_6787; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7824 = _T_5 ? tag_90 : _GEN_6788; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7825 = _T_5 ? tag_91 : _GEN_6789; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7826 = _T_5 ? tag_92 : _GEN_6790; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7827 = _T_5 ? tag_93 : _GEN_6791; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7828 = _T_5 ? tag_94 : _GEN_6792; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7829 = _T_5 ? tag_95 : _GEN_6793; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7830 = _T_5 ? tag_96 : _GEN_6794; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7831 = _T_5 ? tag_97 : _GEN_6795; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7832 = _T_5 ? tag_98 : _GEN_6796; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7833 = _T_5 ? tag_99 : _GEN_6797; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7834 = _T_5 ? tag_100 : _GEN_6798; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7835 = _T_5 ? tag_101 : _GEN_6799; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7836 = _T_5 ? tag_102 : _GEN_6800; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7837 = _T_5 ? tag_103 : _GEN_6801; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7838 = _T_5 ? tag_104 : _GEN_6802; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7839 = _T_5 ? tag_105 : _GEN_6803; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7840 = _T_5 ? tag_106 : _GEN_6804; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7841 = _T_5 ? tag_107 : _GEN_6805; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7842 = _T_5 ? tag_108 : _GEN_6806; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7843 = _T_5 ? tag_109 : _GEN_6807; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7844 = _T_5 ? tag_110 : _GEN_6808; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7845 = _T_5 ? tag_111 : _GEN_6809; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7846 = _T_5 ? tag_112 : _GEN_6810; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7847 = _T_5 ? tag_113 : _GEN_6811; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7848 = _T_5 ? tag_114 : _GEN_6812; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7849 = _T_5 ? tag_115 : _GEN_6813; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7850 = _T_5 ? tag_116 : _GEN_6814; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7851 = _T_5 ? tag_117 : _GEN_6815; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7852 = _T_5 ? tag_118 : _GEN_6816; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7853 = _T_5 ? tag_119 : _GEN_6817; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7854 = _T_5 ? tag_120 : _GEN_6818; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7855 = _T_5 ? tag_121 : _GEN_6819; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7856 = _T_5 ? tag_122 : _GEN_6820; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7857 = _T_5 ? tag_123 : _GEN_6821; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7858 = _T_5 ? tag_124 : _GEN_6822; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7859 = _T_5 ? tag_125 : _GEN_6823; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7860 = _T_5 ? tag_126 : _GEN_6824; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7861 = _T_5 ? tag_127 : _GEN_6825; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7862 = _T_5 ? tag_128 : _GEN_6826; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7863 = _T_5 ? tag_129 : _GEN_6827; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7864 = _T_5 ? tag_130 : _GEN_6828; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7865 = _T_5 ? tag_131 : _GEN_6829; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7866 = _T_5 ? tag_132 : _GEN_6830; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7867 = _T_5 ? tag_133 : _GEN_6831; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7868 = _T_5 ? tag_134 : _GEN_6832; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7869 = _T_5 ? tag_135 : _GEN_6833; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7870 = _T_5 ? tag_136 : _GEN_6834; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7871 = _T_5 ? tag_137 : _GEN_6835; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7872 = _T_5 ? tag_138 : _GEN_6836; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7873 = _T_5 ? tag_139 : _GEN_6837; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7874 = _T_5 ? tag_140 : _GEN_6838; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7875 = _T_5 ? tag_141 : _GEN_6839; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7876 = _T_5 ? tag_142 : _GEN_6840; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7877 = _T_5 ? tag_143 : _GEN_6841; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7878 = _T_5 ? tag_144 : _GEN_6842; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7879 = _T_5 ? tag_145 : _GEN_6843; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7880 = _T_5 ? tag_146 : _GEN_6844; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7881 = _T_5 ? tag_147 : _GEN_6845; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7882 = _T_5 ? tag_148 : _GEN_6846; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7883 = _T_5 ? tag_149 : _GEN_6847; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7884 = _T_5 ? tag_150 : _GEN_6848; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7885 = _T_5 ? tag_151 : _GEN_6849; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7886 = _T_5 ? tag_152 : _GEN_6850; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7887 = _T_5 ? tag_153 : _GEN_6851; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7888 = _T_5 ? tag_154 : _GEN_6852; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7889 = _T_5 ? tag_155 : _GEN_6853; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7890 = _T_5 ? tag_156 : _GEN_6854; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7891 = _T_5 ? tag_157 : _GEN_6855; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7892 = _T_5 ? tag_158 : _GEN_6856; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7893 = _T_5 ? tag_159 : _GEN_6857; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7894 = _T_5 ? tag_160 : _GEN_6858; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7895 = _T_5 ? tag_161 : _GEN_6859; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7896 = _T_5 ? tag_162 : _GEN_6860; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7897 = _T_5 ? tag_163 : _GEN_6861; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7898 = _T_5 ? tag_164 : _GEN_6862; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7899 = _T_5 ? tag_165 : _GEN_6863; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7900 = _T_5 ? tag_166 : _GEN_6864; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7901 = _T_5 ? tag_167 : _GEN_6865; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7902 = _T_5 ? tag_168 : _GEN_6866; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7903 = _T_5 ? tag_169 : _GEN_6867; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7904 = _T_5 ? tag_170 : _GEN_6868; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7905 = _T_5 ? tag_171 : _GEN_6869; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7906 = _T_5 ? tag_172 : _GEN_6870; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7907 = _T_5 ? tag_173 : _GEN_6871; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7908 = _T_5 ? tag_174 : _GEN_6872; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7909 = _T_5 ? tag_175 : _GEN_6873; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7910 = _T_5 ? tag_176 : _GEN_6874; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7911 = _T_5 ? tag_177 : _GEN_6875; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7912 = _T_5 ? tag_178 : _GEN_6876; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7913 = _T_5 ? tag_179 : _GEN_6877; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7914 = _T_5 ? tag_180 : _GEN_6878; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7915 = _T_5 ? tag_181 : _GEN_6879; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7916 = _T_5 ? tag_182 : _GEN_6880; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7917 = _T_5 ? tag_183 : _GEN_6881; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7918 = _T_5 ? tag_184 : _GEN_6882; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7919 = _T_5 ? tag_185 : _GEN_6883; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7920 = _T_5 ? tag_186 : _GEN_6884; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7921 = _T_5 ? tag_187 : _GEN_6885; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7922 = _T_5 ? tag_188 : _GEN_6886; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7923 = _T_5 ? tag_189 : _GEN_6887; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7924 = _T_5 ? tag_190 : _GEN_6888; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7925 = _T_5 ? tag_191 : _GEN_6889; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7926 = _T_5 ? tag_192 : _GEN_6890; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7927 = _T_5 ? tag_193 : _GEN_6891; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7928 = _T_5 ? tag_194 : _GEN_6892; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7929 = _T_5 ? tag_195 : _GEN_6893; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7930 = _T_5 ? tag_196 : _GEN_6894; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7931 = _T_5 ? tag_197 : _GEN_6895; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7932 = _T_5 ? tag_198 : _GEN_6896; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7933 = _T_5 ? tag_199 : _GEN_6897; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7934 = _T_5 ? tag_200 : _GEN_6898; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7935 = _T_5 ? tag_201 : _GEN_6899; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7936 = _T_5 ? tag_202 : _GEN_6900; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7937 = _T_5 ? tag_203 : _GEN_6901; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7938 = _T_5 ? tag_204 : _GEN_6902; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7939 = _T_5 ? tag_205 : _GEN_6903; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7940 = _T_5 ? tag_206 : _GEN_6904; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7941 = _T_5 ? tag_207 : _GEN_6905; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7942 = _T_5 ? tag_208 : _GEN_6906; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7943 = _T_5 ? tag_209 : _GEN_6907; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7944 = _T_5 ? tag_210 : _GEN_6908; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7945 = _T_5 ? tag_211 : _GEN_6909; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7946 = _T_5 ? tag_212 : _GEN_6910; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7947 = _T_5 ? tag_213 : _GEN_6911; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7948 = _T_5 ? tag_214 : _GEN_6912; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7949 = _T_5 ? tag_215 : _GEN_6913; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7950 = _T_5 ? tag_216 : _GEN_6914; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7951 = _T_5 ? tag_217 : _GEN_6915; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7952 = _T_5 ? tag_218 : _GEN_6916; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7953 = _T_5 ? tag_219 : _GEN_6917; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7954 = _T_5 ? tag_220 : _GEN_6918; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7955 = _T_5 ? tag_221 : _GEN_6919; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7956 = _T_5 ? tag_222 : _GEN_6920; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7957 = _T_5 ? tag_223 : _GEN_6921; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7958 = _T_5 ? tag_224 : _GEN_6922; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7959 = _T_5 ? tag_225 : _GEN_6923; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7960 = _T_5 ? tag_226 : _GEN_6924; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7961 = _T_5 ? tag_227 : _GEN_6925; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7962 = _T_5 ? tag_228 : _GEN_6926; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7963 = _T_5 ? tag_229 : _GEN_6927; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7964 = _T_5 ? tag_230 : _GEN_6928; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7965 = _T_5 ? tag_231 : _GEN_6929; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7966 = _T_5 ? tag_232 : _GEN_6930; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7967 = _T_5 ? tag_233 : _GEN_6931; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7968 = _T_5 ? tag_234 : _GEN_6932; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7969 = _T_5 ? tag_235 : _GEN_6933; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7970 = _T_5 ? tag_236 : _GEN_6934; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7971 = _T_5 ? tag_237 : _GEN_6935; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7972 = _T_5 ? tag_238 : _GEN_6936; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7973 = _T_5 ? tag_239 : _GEN_6937; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7974 = _T_5 ? tag_240 : _GEN_6938; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7975 = _T_5 ? tag_241 : _GEN_6939; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7976 = _T_5 ? tag_242 : _GEN_6940; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7977 = _T_5 ? tag_243 : _GEN_6941; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7978 = _T_5 ? tag_244 : _GEN_6942; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7979 = _T_5 ? tag_245 : _GEN_6943; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7980 = _T_5 ? tag_246 : _GEN_6944; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7981 = _T_5 ? tag_247 : _GEN_6945; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7982 = _T_5 ? tag_248 : _GEN_6946; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7983 = _T_5 ? tag_249 : _GEN_6947; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7984 = _T_5 ? tag_250 : _GEN_6948; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7985 = _T_5 ? tag_251 : _GEN_6949; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7986 = _T_5 ? tag_252 : _GEN_6950; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7987 = _T_5 ? tag_253 : _GEN_6951; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7988 = _T_5 ? tag_254 : _GEN_6952; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_7989 = _T_5 ? tag_255 : _GEN_6953; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire  _GEN_7990 = _T_5 ? dirty_0 : _GEN_6954; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7991 = _T_5 ? dirty_1 : _GEN_6955; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7992 = _T_5 ? dirty_2 : _GEN_6956; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7993 = _T_5 ? dirty_3 : _GEN_6957; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7994 = _T_5 ? dirty_4 : _GEN_6958; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7995 = _T_5 ? dirty_5 : _GEN_6959; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7996 = _T_5 ? dirty_6 : _GEN_6960; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7997 = _T_5 ? dirty_7 : _GEN_6961; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7998 = _T_5 ? dirty_8 : _GEN_6962; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7999 = _T_5 ? dirty_9 : _GEN_6963; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8000 = _T_5 ? dirty_10 : _GEN_6964; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8001 = _T_5 ? dirty_11 : _GEN_6965; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8002 = _T_5 ? dirty_12 : _GEN_6966; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8003 = _T_5 ? dirty_13 : _GEN_6967; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8004 = _T_5 ? dirty_14 : _GEN_6968; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8005 = _T_5 ? dirty_15 : _GEN_6969; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8006 = _T_5 ? dirty_16 : _GEN_6970; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8007 = _T_5 ? dirty_17 : _GEN_6971; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8008 = _T_5 ? dirty_18 : _GEN_6972; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8009 = _T_5 ? dirty_19 : _GEN_6973; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8010 = _T_5 ? dirty_20 : _GEN_6974; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8011 = _T_5 ? dirty_21 : _GEN_6975; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8012 = _T_5 ? dirty_22 : _GEN_6976; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8013 = _T_5 ? dirty_23 : _GEN_6977; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8014 = _T_5 ? dirty_24 : _GEN_6978; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8015 = _T_5 ? dirty_25 : _GEN_6979; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8016 = _T_5 ? dirty_26 : _GEN_6980; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8017 = _T_5 ? dirty_27 : _GEN_6981; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8018 = _T_5 ? dirty_28 : _GEN_6982; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8019 = _T_5 ? dirty_29 : _GEN_6983; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8020 = _T_5 ? dirty_30 : _GEN_6984; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8021 = _T_5 ? dirty_31 : _GEN_6985; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8022 = _T_5 ? dirty_32 : _GEN_6986; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8023 = _T_5 ? dirty_33 : _GEN_6987; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8024 = _T_5 ? dirty_34 : _GEN_6988; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8025 = _T_5 ? dirty_35 : _GEN_6989; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8026 = _T_5 ? dirty_36 : _GEN_6990; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8027 = _T_5 ? dirty_37 : _GEN_6991; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8028 = _T_5 ? dirty_38 : _GEN_6992; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8029 = _T_5 ? dirty_39 : _GEN_6993; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8030 = _T_5 ? dirty_40 : _GEN_6994; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8031 = _T_5 ? dirty_41 : _GEN_6995; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8032 = _T_5 ? dirty_42 : _GEN_6996; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8033 = _T_5 ? dirty_43 : _GEN_6997; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8034 = _T_5 ? dirty_44 : _GEN_6998; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8035 = _T_5 ? dirty_45 : _GEN_6999; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8036 = _T_5 ? dirty_46 : _GEN_7000; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8037 = _T_5 ? dirty_47 : _GEN_7001; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8038 = _T_5 ? dirty_48 : _GEN_7002; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8039 = _T_5 ? dirty_49 : _GEN_7003; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8040 = _T_5 ? dirty_50 : _GEN_7004; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8041 = _T_5 ? dirty_51 : _GEN_7005; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8042 = _T_5 ? dirty_52 : _GEN_7006; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8043 = _T_5 ? dirty_53 : _GEN_7007; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8044 = _T_5 ? dirty_54 : _GEN_7008; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8045 = _T_5 ? dirty_55 : _GEN_7009; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8046 = _T_5 ? dirty_56 : _GEN_7010; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8047 = _T_5 ? dirty_57 : _GEN_7011; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8048 = _T_5 ? dirty_58 : _GEN_7012; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8049 = _T_5 ? dirty_59 : _GEN_7013; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8050 = _T_5 ? dirty_60 : _GEN_7014; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8051 = _T_5 ? dirty_61 : _GEN_7015; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8052 = _T_5 ? dirty_62 : _GEN_7016; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8053 = _T_5 ? dirty_63 : _GEN_7017; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8054 = _T_5 ? dirty_64 : _GEN_7018; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8055 = _T_5 ? dirty_65 : _GEN_7019; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8056 = _T_5 ? dirty_66 : _GEN_7020; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8057 = _T_5 ? dirty_67 : _GEN_7021; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8058 = _T_5 ? dirty_68 : _GEN_7022; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8059 = _T_5 ? dirty_69 : _GEN_7023; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8060 = _T_5 ? dirty_70 : _GEN_7024; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8061 = _T_5 ? dirty_71 : _GEN_7025; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8062 = _T_5 ? dirty_72 : _GEN_7026; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8063 = _T_5 ? dirty_73 : _GEN_7027; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8064 = _T_5 ? dirty_74 : _GEN_7028; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8065 = _T_5 ? dirty_75 : _GEN_7029; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8066 = _T_5 ? dirty_76 : _GEN_7030; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8067 = _T_5 ? dirty_77 : _GEN_7031; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8068 = _T_5 ? dirty_78 : _GEN_7032; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8069 = _T_5 ? dirty_79 : _GEN_7033; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8070 = _T_5 ? dirty_80 : _GEN_7034; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8071 = _T_5 ? dirty_81 : _GEN_7035; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8072 = _T_5 ? dirty_82 : _GEN_7036; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8073 = _T_5 ? dirty_83 : _GEN_7037; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8074 = _T_5 ? dirty_84 : _GEN_7038; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8075 = _T_5 ? dirty_85 : _GEN_7039; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8076 = _T_5 ? dirty_86 : _GEN_7040; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8077 = _T_5 ? dirty_87 : _GEN_7041; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8078 = _T_5 ? dirty_88 : _GEN_7042; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8079 = _T_5 ? dirty_89 : _GEN_7043; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8080 = _T_5 ? dirty_90 : _GEN_7044; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8081 = _T_5 ? dirty_91 : _GEN_7045; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8082 = _T_5 ? dirty_92 : _GEN_7046; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8083 = _T_5 ? dirty_93 : _GEN_7047; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8084 = _T_5 ? dirty_94 : _GEN_7048; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8085 = _T_5 ? dirty_95 : _GEN_7049; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8086 = _T_5 ? dirty_96 : _GEN_7050; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8087 = _T_5 ? dirty_97 : _GEN_7051; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8088 = _T_5 ? dirty_98 : _GEN_7052; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8089 = _T_5 ? dirty_99 : _GEN_7053; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8090 = _T_5 ? dirty_100 : _GEN_7054; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8091 = _T_5 ? dirty_101 : _GEN_7055; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8092 = _T_5 ? dirty_102 : _GEN_7056; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8093 = _T_5 ? dirty_103 : _GEN_7057; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8094 = _T_5 ? dirty_104 : _GEN_7058; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8095 = _T_5 ? dirty_105 : _GEN_7059; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8096 = _T_5 ? dirty_106 : _GEN_7060; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8097 = _T_5 ? dirty_107 : _GEN_7061; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8098 = _T_5 ? dirty_108 : _GEN_7062; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8099 = _T_5 ? dirty_109 : _GEN_7063; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8100 = _T_5 ? dirty_110 : _GEN_7064; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8101 = _T_5 ? dirty_111 : _GEN_7065; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8102 = _T_5 ? dirty_112 : _GEN_7066; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8103 = _T_5 ? dirty_113 : _GEN_7067; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8104 = _T_5 ? dirty_114 : _GEN_7068; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8105 = _T_5 ? dirty_115 : _GEN_7069; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8106 = _T_5 ? dirty_116 : _GEN_7070; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8107 = _T_5 ? dirty_117 : _GEN_7071; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8108 = _T_5 ? dirty_118 : _GEN_7072; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8109 = _T_5 ? dirty_119 : _GEN_7073; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8110 = _T_5 ? dirty_120 : _GEN_7074; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8111 = _T_5 ? dirty_121 : _GEN_7075; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8112 = _T_5 ? dirty_122 : _GEN_7076; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8113 = _T_5 ? dirty_123 : _GEN_7077; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8114 = _T_5 ? dirty_124 : _GEN_7078; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8115 = _T_5 ? dirty_125 : _GEN_7079; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8116 = _T_5 ? dirty_126 : _GEN_7080; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8117 = _T_5 ? dirty_127 : _GEN_7081; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8118 = _T_5 ? dirty_128 : _GEN_7082; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8119 = _T_5 ? dirty_129 : _GEN_7083; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8120 = _T_5 ? dirty_130 : _GEN_7084; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8121 = _T_5 ? dirty_131 : _GEN_7085; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8122 = _T_5 ? dirty_132 : _GEN_7086; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8123 = _T_5 ? dirty_133 : _GEN_7087; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8124 = _T_5 ? dirty_134 : _GEN_7088; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8125 = _T_5 ? dirty_135 : _GEN_7089; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8126 = _T_5 ? dirty_136 : _GEN_7090; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8127 = _T_5 ? dirty_137 : _GEN_7091; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8128 = _T_5 ? dirty_138 : _GEN_7092; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8129 = _T_5 ? dirty_139 : _GEN_7093; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8130 = _T_5 ? dirty_140 : _GEN_7094; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8131 = _T_5 ? dirty_141 : _GEN_7095; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8132 = _T_5 ? dirty_142 : _GEN_7096; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8133 = _T_5 ? dirty_143 : _GEN_7097; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8134 = _T_5 ? dirty_144 : _GEN_7098; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8135 = _T_5 ? dirty_145 : _GEN_7099; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8136 = _T_5 ? dirty_146 : _GEN_7100; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8137 = _T_5 ? dirty_147 : _GEN_7101; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8138 = _T_5 ? dirty_148 : _GEN_7102; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8139 = _T_5 ? dirty_149 : _GEN_7103; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8140 = _T_5 ? dirty_150 : _GEN_7104; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8141 = _T_5 ? dirty_151 : _GEN_7105; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8142 = _T_5 ? dirty_152 : _GEN_7106; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8143 = _T_5 ? dirty_153 : _GEN_7107; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8144 = _T_5 ? dirty_154 : _GEN_7108; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8145 = _T_5 ? dirty_155 : _GEN_7109; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8146 = _T_5 ? dirty_156 : _GEN_7110; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8147 = _T_5 ? dirty_157 : _GEN_7111; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8148 = _T_5 ? dirty_158 : _GEN_7112; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8149 = _T_5 ? dirty_159 : _GEN_7113; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8150 = _T_5 ? dirty_160 : _GEN_7114; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8151 = _T_5 ? dirty_161 : _GEN_7115; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8152 = _T_5 ? dirty_162 : _GEN_7116; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8153 = _T_5 ? dirty_163 : _GEN_7117; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8154 = _T_5 ? dirty_164 : _GEN_7118; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8155 = _T_5 ? dirty_165 : _GEN_7119; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8156 = _T_5 ? dirty_166 : _GEN_7120; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8157 = _T_5 ? dirty_167 : _GEN_7121; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8158 = _T_5 ? dirty_168 : _GEN_7122; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8159 = _T_5 ? dirty_169 : _GEN_7123; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8160 = _T_5 ? dirty_170 : _GEN_7124; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8161 = _T_5 ? dirty_171 : _GEN_7125; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8162 = _T_5 ? dirty_172 : _GEN_7126; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8163 = _T_5 ? dirty_173 : _GEN_7127; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8164 = _T_5 ? dirty_174 : _GEN_7128; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8165 = _T_5 ? dirty_175 : _GEN_7129; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8166 = _T_5 ? dirty_176 : _GEN_7130; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8167 = _T_5 ? dirty_177 : _GEN_7131; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8168 = _T_5 ? dirty_178 : _GEN_7132; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8169 = _T_5 ? dirty_179 : _GEN_7133; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8170 = _T_5 ? dirty_180 : _GEN_7134; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8171 = _T_5 ? dirty_181 : _GEN_7135; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8172 = _T_5 ? dirty_182 : _GEN_7136; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8173 = _T_5 ? dirty_183 : _GEN_7137; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8174 = _T_5 ? dirty_184 : _GEN_7138; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8175 = _T_5 ? dirty_185 : _GEN_7139; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8176 = _T_5 ? dirty_186 : _GEN_7140; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8177 = _T_5 ? dirty_187 : _GEN_7141; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8178 = _T_5 ? dirty_188 : _GEN_7142; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8179 = _T_5 ? dirty_189 : _GEN_7143; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8180 = _T_5 ? dirty_190 : _GEN_7144; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8181 = _T_5 ? dirty_191 : _GEN_7145; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8182 = _T_5 ? dirty_192 : _GEN_7146; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8183 = _T_5 ? dirty_193 : _GEN_7147; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8184 = _T_5 ? dirty_194 : _GEN_7148; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8185 = _T_5 ? dirty_195 : _GEN_7149; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8186 = _T_5 ? dirty_196 : _GEN_7150; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8187 = _T_5 ? dirty_197 : _GEN_7151; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8188 = _T_5 ? dirty_198 : _GEN_7152; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8189 = _T_5 ? dirty_199 : _GEN_7153; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8190 = _T_5 ? dirty_200 : _GEN_7154; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8191 = _T_5 ? dirty_201 : _GEN_7155; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8192 = _T_5 ? dirty_202 : _GEN_7156; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8193 = _T_5 ? dirty_203 : _GEN_7157; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8194 = _T_5 ? dirty_204 : _GEN_7158; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8195 = _T_5 ? dirty_205 : _GEN_7159; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8196 = _T_5 ? dirty_206 : _GEN_7160; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8197 = _T_5 ? dirty_207 : _GEN_7161; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8198 = _T_5 ? dirty_208 : _GEN_7162; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8199 = _T_5 ? dirty_209 : _GEN_7163; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8200 = _T_5 ? dirty_210 : _GEN_7164; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8201 = _T_5 ? dirty_211 : _GEN_7165; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8202 = _T_5 ? dirty_212 : _GEN_7166; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8203 = _T_5 ? dirty_213 : _GEN_7167; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8204 = _T_5 ? dirty_214 : _GEN_7168; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8205 = _T_5 ? dirty_215 : _GEN_7169; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8206 = _T_5 ? dirty_216 : _GEN_7170; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8207 = _T_5 ? dirty_217 : _GEN_7171; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8208 = _T_5 ? dirty_218 : _GEN_7172; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8209 = _T_5 ? dirty_219 : _GEN_7173; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8210 = _T_5 ? dirty_220 : _GEN_7174; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8211 = _T_5 ? dirty_221 : _GEN_7175; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8212 = _T_5 ? dirty_222 : _GEN_7176; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8213 = _T_5 ? dirty_223 : _GEN_7177; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8214 = _T_5 ? dirty_224 : _GEN_7178; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8215 = _T_5 ? dirty_225 : _GEN_7179; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8216 = _T_5 ? dirty_226 : _GEN_7180; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8217 = _T_5 ? dirty_227 : _GEN_7181; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8218 = _T_5 ? dirty_228 : _GEN_7182; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8219 = _T_5 ? dirty_229 : _GEN_7183; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8220 = _T_5 ? dirty_230 : _GEN_7184; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8221 = _T_5 ? dirty_231 : _GEN_7185; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8222 = _T_5 ? dirty_232 : _GEN_7186; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8223 = _T_5 ? dirty_233 : _GEN_7187; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8224 = _T_5 ? dirty_234 : _GEN_7188; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8225 = _T_5 ? dirty_235 : _GEN_7189; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8226 = _T_5 ? dirty_236 : _GEN_7190; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8227 = _T_5 ? dirty_237 : _GEN_7191; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8228 = _T_5 ? dirty_238 : _GEN_7192; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8229 = _T_5 ? dirty_239 : _GEN_7193; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8230 = _T_5 ? dirty_240 : _GEN_7194; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8231 = _T_5 ? dirty_241 : _GEN_7195; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8232 = _T_5 ? dirty_242 : _GEN_7196; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8233 = _T_5 ? dirty_243 : _GEN_7197; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8234 = _T_5 ? dirty_244 : _GEN_7198; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8235 = _T_5 ? dirty_245 : _GEN_7199; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8236 = _T_5 ? dirty_246 : _GEN_7200; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8237 = _T_5 ? dirty_247 : _GEN_7201; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8238 = _T_5 ? dirty_248 : _GEN_7202; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8239 = _T_5 ? dirty_249 : _GEN_7203; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8240 = _T_5 ? dirty_250 : _GEN_7204; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8241 = _T_5 ? dirty_251 : _GEN_7205; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8242 = _T_5 ? dirty_252 : _GEN_7206; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8243 = _T_5 ? dirty_253 : _GEN_7207; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8244 = _T_5 ? dirty_254 : _GEN_7208; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_8245 = _T_5 ? dirty_255 : _GEN_7209; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire [3:0] _GEN_8246 = _T_5 ? offset_0 : _GEN_7210; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8247 = _T_5 ? offset_1 : _GEN_7211; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8248 = _T_5 ? offset_2 : _GEN_7212; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8249 = _T_5 ? offset_3 : _GEN_7213; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8250 = _T_5 ? offset_4 : _GEN_7214; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8251 = _T_5 ? offset_5 : _GEN_7215; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8252 = _T_5 ? offset_6 : _GEN_7216; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8253 = _T_5 ? offset_7 : _GEN_7217; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8254 = _T_5 ? offset_8 : _GEN_7218; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8255 = _T_5 ? offset_9 : _GEN_7219; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8256 = _T_5 ? offset_10 : _GEN_7220; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8257 = _T_5 ? offset_11 : _GEN_7221; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8258 = _T_5 ? offset_12 : _GEN_7222; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8259 = _T_5 ? offset_13 : _GEN_7223; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8260 = _T_5 ? offset_14 : _GEN_7224; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8261 = _T_5 ? offset_15 : _GEN_7225; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8262 = _T_5 ? offset_16 : _GEN_7226; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8263 = _T_5 ? offset_17 : _GEN_7227; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8264 = _T_5 ? offset_18 : _GEN_7228; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8265 = _T_5 ? offset_19 : _GEN_7229; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8266 = _T_5 ? offset_20 : _GEN_7230; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8267 = _T_5 ? offset_21 : _GEN_7231; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8268 = _T_5 ? offset_22 : _GEN_7232; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8269 = _T_5 ? offset_23 : _GEN_7233; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8270 = _T_5 ? offset_24 : _GEN_7234; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8271 = _T_5 ? offset_25 : _GEN_7235; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8272 = _T_5 ? offset_26 : _GEN_7236; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8273 = _T_5 ? offset_27 : _GEN_7237; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8274 = _T_5 ? offset_28 : _GEN_7238; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8275 = _T_5 ? offset_29 : _GEN_7239; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8276 = _T_5 ? offset_30 : _GEN_7240; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8277 = _T_5 ? offset_31 : _GEN_7241; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8278 = _T_5 ? offset_32 : _GEN_7242; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8279 = _T_5 ? offset_33 : _GEN_7243; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8280 = _T_5 ? offset_34 : _GEN_7244; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8281 = _T_5 ? offset_35 : _GEN_7245; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8282 = _T_5 ? offset_36 : _GEN_7246; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8283 = _T_5 ? offset_37 : _GEN_7247; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8284 = _T_5 ? offset_38 : _GEN_7248; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8285 = _T_5 ? offset_39 : _GEN_7249; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8286 = _T_5 ? offset_40 : _GEN_7250; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8287 = _T_5 ? offset_41 : _GEN_7251; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8288 = _T_5 ? offset_42 : _GEN_7252; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8289 = _T_5 ? offset_43 : _GEN_7253; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8290 = _T_5 ? offset_44 : _GEN_7254; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8291 = _T_5 ? offset_45 : _GEN_7255; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8292 = _T_5 ? offset_46 : _GEN_7256; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8293 = _T_5 ? offset_47 : _GEN_7257; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8294 = _T_5 ? offset_48 : _GEN_7258; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8295 = _T_5 ? offset_49 : _GEN_7259; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8296 = _T_5 ? offset_50 : _GEN_7260; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8297 = _T_5 ? offset_51 : _GEN_7261; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8298 = _T_5 ? offset_52 : _GEN_7262; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8299 = _T_5 ? offset_53 : _GEN_7263; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8300 = _T_5 ? offset_54 : _GEN_7264; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8301 = _T_5 ? offset_55 : _GEN_7265; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8302 = _T_5 ? offset_56 : _GEN_7266; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8303 = _T_5 ? offset_57 : _GEN_7267; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8304 = _T_5 ? offset_58 : _GEN_7268; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8305 = _T_5 ? offset_59 : _GEN_7269; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8306 = _T_5 ? offset_60 : _GEN_7270; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8307 = _T_5 ? offset_61 : _GEN_7271; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8308 = _T_5 ? offset_62 : _GEN_7272; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8309 = _T_5 ? offset_63 : _GEN_7273; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8310 = _T_5 ? offset_64 : _GEN_7274; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8311 = _T_5 ? offset_65 : _GEN_7275; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8312 = _T_5 ? offset_66 : _GEN_7276; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8313 = _T_5 ? offset_67 : _GEN_7277; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8314 = _T_5 ? offset_68 : _GEN_7278; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8315 = _T_5 ? offset_69 : _GEN_7279; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8316 = _T_5 ? offset_70 : _GEN_7280; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8317 = _T_5 ? offset_71 : _GEN_7281; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8318 = _T_5 ? offset_72 : _GEN_7282; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8319 = _T_5 ? offset_73 : _GEN_7283; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8320 = _T_5 ? offset_74 : _GEN_7284; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8321 = _T_5 ? offset_75 : _GEN_7285; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8322 = _T_5 ? offset_76 : _GEN_7286; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8323 = _T_5 ? offset_77 : _GEN_7287; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8324 = _T_5 ? offset_78 : _GEN_7288; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8325 = _T_5 ? offset_79 : _GEN_7289; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8326 = _T_5 ? offset_80 : _GEN_7290; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8327 = _T_5 ? offset_81 : _GEN_7291; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8328 = _T_5 ? offset_82 : _GEN_7292; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8329 = _T_5 ? offset_83 : _GEN_7293; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8330 = _T_5 ? offset_84 : _GEN_7294; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8331 = _T_5 ? offset_85 : _GEN_7295; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8332 = _T_5 ? offset_86 : _GEN_7296; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8333 = _T_5 ? offset_87 : _GEN_7297; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8334 = _T_5 ? offset_88 : _GEN_7298; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8335 = _T_5 ? offset_89 : _GEN_7299; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8336 = _T_5 ? offset_90 : _GEN_7300; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8337 = _T_5 ? offset_91 : _GEN_7301; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8338 = _T_5 ? offset_92 : _GEN_7302; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8339 = _T_5 ? offset_93 : _GEN_7303; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8340 = _T_5 ? offset_94 : _GEN_7304; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8341 = _T_5 ? offset_95 : _GEN_7305; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8342 = _T_5 ? offset_96 : _GEN_7306; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8343 = _T_5 ? offset_97 : _GEN_7307; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8344 = _T_5 ? offset_98 : _GEN_7308; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8345 = _T_5 ? offset_99 : _GEN_7309; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8346 = _T_5 ? offset_100 : _GEN_7310; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8347 = _T_5 ? offset_101 : _GEN_7311; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8348 = _T_5 ? offset_102 : _GEN_7312; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8349 = _T_5 ? offset_103 : _GEN_7313; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8350 = _T_5 ? offset_104 : _GEN_7314; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8351 = _T_5 ? offset_105 : _GEN_7315; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8352 = _T_5 ? offset_106 : _GEN_7316; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8353 = _T_5 ? offset_107 : _GEN_7317; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8354 = _T_5 ? offset_108 : _GEN_7318; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8355 = _T_5 ? offset_109 : _GEN_7319; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8356 = _T_5 ? offset_110 : _GEN_7320; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8357 = _T_5 ? offset_111 : _GEN_7321; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8358 = _T_5 ? offset_112 : _GEN_7322; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8359 = _T_5 ? offset_113 : _GEN_7323; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8360 = _T_5 ? offset_114 : _GEN_7324; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8361 = _T_5 ? offset_115 : _GEN_7325; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8362 = _T_5 ? offset_116 : _GEN_7326; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8363 = _T_5 ? offset_117 : _GEN_7327; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8364 = _T_5 ? offset_118 : _GEN_7328; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8365 = _T_5 ? offset_119 : _GEN_7329; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8366 = _T_5 ? offset_120 : _GEN_7330; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8367 = _T_5 ? offset_121 : _GEN_7331; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8368 = _T_5 ? offset_122 : _GEN_7332; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8369 = _T_5 ? offset_123 : _GEN_7333; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8370 = _T_5 ? offset_124 : _GEN_7334; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8371 = _T_5 ? offset_125 : _GEN_7335; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8372 = _T_5 ? offset_126 : _GEN_7336; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8373 = _T_5 ? offset_127 : _GEN_7337; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8374 = _T_5 ? offset_128 : _GEN_7338; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8375 = _T_5 ? offset_129 : _GEN_7339; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8376 = _T_5 ? offset_130 : _GEN_7340; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8377 = _T_5 ? offset_131 : _GEN_7341; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8378 = _T_5 ? offset_132 : _GEN_7342; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8379 = _T_5 ? offset_133 : _GEN_7343; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8380 = _T_5 ? offset_134 : _GEN_7344; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8381 = _T_5 ? offset_135 : _GEN_7345; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8382 = _T_5 ? offset_136 : _GEN_7346; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8383 = _T_5 ? offset_137 : _GEN_7347; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8384 = _T_5 ? offset_138 : _GEN_7348; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8385 = _T_5 ? offset_139 : _GEN_7349; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8386 = _T_5 ? offset_140 : _GEN_7350; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8387 = _T_5 ? offset_141 : _GEN_7351; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8388 = _T_5 ? offset_142 : _GEN_7352; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8389 = _T_5 ? offset_143 : _GEN_7353; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8390 = _T_5 ? offset_144 : _GEN_7354; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8391 = _T_5 ? offset_145 : _GEN_7355; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8392 = _T_5 ? offset_146 : _GEN_7356; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8393 = _T_5 ? offset_147 : _GEN_7357; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8394 = _T_5 ? offset_148 : _GEN_7358; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8395 = _T_5 ? offset_149 : _GEN_7359; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8396 = _T_5 ? offset_150 : _GEN_7360; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8397 = _T_5 ? offset_151 : _GEN_7361; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8398 = _T_5 ? offset_152 : _GEN_7362; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8399 = _T_5 ? offset_153 : _GEN_7363; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8400 = _T_5 ? offset_154 : _GEN_7364; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8401 = _T_5 ? offset_155 : _GEN_7365; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8402 = _T_5 ? offset_156 : _GEN_7366; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8403 = _T_5 ? offset_157 : _GEN_7367; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8404 = _T_5 ? offset_158 : _GEN_7368; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8405 = _T_5 ? offset_159 : _GEN_7369; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8406 = _T_5 ? offset_160 : _GEN_7370; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8407 = _T_5 ? offset_161 : _GEN_7371; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8408 = _T_5 ? offset_162 : _GEN_7372; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8409 = _T_5 ? offset_163 : _GEN_7373; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8410 = _T_5 ? offset_164 : _GEN_7374; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8411 = _T_5 ? offset_165 : _GEN_7375; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8412 = _T_5 ? offset_166 : _GEN_7376; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8413 = _T_5 ? offset_167 : _GEN_7377; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8414 = _T_5 ? offset_168 : _GEN_7378; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8415 = _T_5 ? offset_169 : _GEN_7379; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8416 = _T_5 ? offset_170 : _GEN_7380; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8417 = _T_5 ? offset_171 : _GEN_7381; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8418 = _T_5 ? offset_172 : _GEN_7382; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8419 = _T_5 ? offset_173 : _GEN_7383; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8420 = _T_5 ? offset_174 : _GEN_7384; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8421 = _T_5 ? offset_175 : _GEN_7385; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8422 = _T_5 ? offset_176 : _GEN_7386; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8423 = _T_5 ? offset_177 : _GEN_7387; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8424 = _T_5 ? offset_178 : _GEN_7388; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8425 = _T_5 ? offset_179 : _GEN_7389; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8426 = _T_5 ? offset_180 : _GEN_7390; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8427 = _T_5 ? offset_181 : _GEN_7391; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8428 = _T_5 ? offset_182 : _GEN_7392; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8429 = _T_5 ? offset_183 : _GEN_7393; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8430 = _T_5 ? offset_184 : _GEN_7394; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8431 = _T_5 ? offset_185 : _GEN_7395; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8432 = _T_5 ? offset_186 : _GEN_7396; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8433 = _T_5 ? offset_187 : _GEN_7397; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8434 = _T_5 ? offset_188 : _GEN_7398; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8435 = _T_5 ? offset_189 : _GEN_7399; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8436 = _T_5 ? offset_190 : _GEN_7400; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8437 = _T_5 ? offset_191 : _GEN_7401; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8438 = _T_5 ? offset_192 : _GEN_7402; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8439 = _T_5 ? offset_193 : _GEN_7403; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8440 = _T_5 ? offset_194 : _GEN_7404; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8441 = _T_5 ? offset_195 : _GEN_7405; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8442 = _T_5 ? offset_196 : _GEN_7406; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8443 = _T_5 ? offset_197 : _GEN_7407; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8444 = _T_5 ? offset_198 : _GEN_7408; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8445 = _T_5 ? offset_199 : _GEN_7409; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8446 = _T_5 ? offset_200 : _GEN_7410; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8447 = _T_5 ? offset_201 : _GEN_7411; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8448 = _T_5 ? offset_202 : _GEN_7412; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8449 = _T_5 ? offset_203 : _GEN_7413; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8450 = _T_5 ? offset_204 : _GEN_7414; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8451 = _T_5 ? offset_205 : _GEN_7415; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8452 = _T_5 ? offset_206 : _GEN_7416; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8453 = _T_5 ? offset_207 : _GEN_7417; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8454 = _T_5 ? offset_208 : _GEN_7418; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8455 = _T_5 ? offset_209 : _GEN_7419; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8456 = _T_5 ? offset_210 : _GEN_7420; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8457 = _T_5 ? offset_211 : _GEN_7421; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8458 = _T_5 ? offset_212 : _GEN_7422; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8459 = _T_5 ? offset_213 : _GEN_7423; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8460 = _T_5 ? offset_214 : _GEN_7424; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8461 = _T_5 ? offset_215 : _GEN_7425; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8462 = _T_5 ? offset_216 : _GEN_7426; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8463 = _T_5 ? offset_217 : _GEN_7427; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8464 = _T_5 ? offset_218 : _GEN_7428; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8465 = _T_5 ? offset_219 : _GEN_7429; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8466 = _T_5 ? offset_220 : _GEN_7430; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8467 = _T_5 ? offset_221 : _GEN_7431; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8468 = _T_5 ? offset_222 : _GEN_7432; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8469 = _T_5 ? offset_223 : _GEN_7433; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8470 = _T_5 ? offset_224 : _GEN_7434; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8471 = _T_5 ? offset_225 : _GEN_7435; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8472 = _T_5 ? offset_226 : _GEN_7436; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8473 = _T_5 ? offset_227 : _GEN_7437; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8474 = _T_5 ? offset_228 : _GEN_7438; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8475 = _T_5 ? offset_229 : _GEN_7439; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8476 = _T_5 ? offset_230 : _GEN_7440; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8477 = _T_5 ? offset_231 : _GEN_7441; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8478 = _T_5 ? offset_232 : _GEN_7442; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8479 = _T_5 ? offset_233 : _GEN_7443; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8480 = _T_5 ? offset_234 : _GEN_7444; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8481 = _T_5 ? offset_235 : _GEN_7445; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8482 = _T_5 ? offset_236 : _GEN_7446; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8483 = _T_5 ? offset_237 : _GEN_7447; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8484 = _T_5 ? offset_238 : _GEN_7448; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8485 = _T_5 ? offset_239 : _GEN_7449; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8486 = _T_5 ? offset_240 : _GEN_7450; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8487 = _T_5 ? offset_241 : _GEN_7451; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8488 = _T_5 ? offset_242 : _GEN_7452; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8489 = _T_5 ? offset_243 : _GEN_7453; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8490 = _T_5 ? offset_244 : _GEN_7454; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8491 = _T_5 ? offset_245 : _GEN_7455; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8492 = _T_5 ? offset_246 : _GEN_7456; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8493 = _T_5 ? offset_247 : _GEN_7457; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8494 = _T_5 ? offset_248 : _GEN_7458; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8495 = _T_5 ? offset_249 : _GEN_7459; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8496 = _T_5 ? offset_250 : _GEN_7460; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8497 = _T_5 ? offset_251 : _GEN_7461; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8498 = _T_5 ? offset_252 : _GEN_7462; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8499 = _T_5 ? offset_253 : _GEN_7463; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8500 = _T_5 ? offset_254 : _GEN_7464; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_8501 = _T_5 ? offset_255 : _GEN_7465; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [31:0] _GEN_8502 = _T_4 ? _data_addr_T : _GEN_7467; // @[Conditional.scala 39:67 Dcache.scala 156:21]
  wire [127:0] _GEN_8503 = _T_4 ? cache_data_out : 128'h0; // @[Conditional.scala 39:67 Dcache.scala 157:21]
  wire [7:0] _GEN_8504 = _T_4 ? 8'hff : 8'h0; // @[Conditional.scala 39:67 Dcache.scala 158:21]
  wire  _GEN_8506 = _T_4 ? _GEN_4365 : _GEN_7471; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_10567 = _T_1 ? 32'h0 : _GEN_8502; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_10568 = _T_1 ? 128'h0 : _GEN_8503; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_10569 = _T_1 ? 8'h0 : _GEN_8504; // @[Conditional.scala 39:67]
  wire  _GEN_10571 = _T_1 ? 1'h0 : _GEN_8506; // @[Conditional.scala 39:67]
  wire  _GEN_10572 = _T_1 ? 1'h0 : _T_4 & _GEN_4365; // @[Conditional.scala 39:67]
  S011HD1P_X32Y2D128_BW req ( // @[Dcache.scala 220:19]
    .Q(req_Q),
    .CLK(req_CLK),
    .CEN(req_CEN),
    .WEN(req_WEN),
    .BWEN(req_BWEN),
    .A(req_A),
    .D(req_D)
  );
  assign io_dmem_data_ready = data_ready; // @[Dcache.scala 217:19]
  assign io_dmem_data_read = 2'h3 == io_dmem_data_size ? valid_rdata : {{31'd0}, _data_read_T_42}; // @[Mux.scala 80:57]
  assign io_out_data_valid = _T ? 1'h0 : _GEN_10571; // @[Conditional.scala 40:58]
  assign io_out_data_req = _T ? 1'h0 : _GEN_10572; // @[Conditional.scala 40:58]
  assign io_out_data_addr = _T ? 32'h0 : _GEN_10567; // @[Conditional.scala 40:58]
  assign io_out_data_strb = _T ? 8'h0 : _GEN_10569; // @[Conditional.scala 40:58]
  assign io_out_data_write = _T ? 128'h0 : _GEN_10568; // @[Conditional.scala 40:58]
  assign req_CLK = clock; // @[Dcache.scala 221:17]
  assign req_CEN = 1'h1; // @[Dcache.scala 222:17]
  assign req_WEN = cache_wen; // @[Dcache.scala 223:17]
  assign req_BWEN = cache_strb; // @[Dcache.scala 224:17]
  assign req_A = io_dmem_data_addr[11:4]; // @[Dcache.scala 29:30]
  assign req_D = cache_wdata; // @[Dcache.scala 226:17]
  always @(posedge clock) begin
    if (reset) begin // @[Dcache.scala 16:24]
      tag_0 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_0 <= _GEN_2306;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_0 <= _GEN_7734;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_1 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_1 <= _GEN_2307;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_1 <= _GEN_7735;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_2 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_2 <= _GEN_2308;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_2 <= _GEN_7736;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_3 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_3 <= _GEN_2309;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_3 <= _GEN_7737;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_4 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_4 <= _GEN_2310;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_4 <= _GEN_7738;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_5 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_5 <= _GEN_2311;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_5 <= _GEN_7739;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_6 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_6 <= _GEN_2312;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_6 <= _GEN_7740;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_7 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_7 <= _GEN_2313;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_7 <= _GEN_7741;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_8 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_8 <= _GEN_2314;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_8 <= _GEN_7742;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_9 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_9 <= _GEN_2315;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_9 <= _GEN_7743;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_10 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_10 <= _GEN_2316;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_10 <= _GEN_7744;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_11 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_11 <= _GEN_2317;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_11 <= _GEN_7745;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_12 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_12 <= _GEN_2318;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_12 <= _GEN_7746;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_13 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_13 <= _GEN_2319;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_13 <= _GEN_7747;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_14 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_14 <= _GEN_2320;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_14 <= _GEN_7748;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_15 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_15 <= _GEN_2321;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_15 <= _GEN_7749;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_16 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_16 <= _GEN_2322;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_16 <= _GEN_7750;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_17 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_17 <= _GEN_2323;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_17 <= _GEN_7751;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_18 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_18 <= _GEN_2324;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_18 <= _GEN_7752;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_19 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_19 <= _GEN_2325;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_19 <= _GEN_7753;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_20 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_20 <= _GEN_2326;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_20 <= _GEN_7754;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_21 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_21 <= _GEN_2327;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_21 <= _GEN_7755;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_22 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_22 <= _GEN_2328;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_22 <= _GEN_7756;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_23 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_23 <= _GEN_2329;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_23 <= _GEN_7757;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_24 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_24 <= _GEN_2330;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_24 <= _GEN_7758;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_25 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_25 <= _GEN_2331;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_25 <= _GEN_7759;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_26 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_26 <= _GEN_2332;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_26 <= _GEN_7760;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_27 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_27 <= _GEN_2333;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_27 <= _GEN_7761;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_28 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_28 <= _GEN_2334;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_28 <= _GEN_7762;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_29 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_29 <= _GEN_2335;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_29 <= _GEN_7763;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_30 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_30 <= _GEN_2336;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_30 <= _GEN_7764;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_31 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_31 <= _GEN_2337;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_31 <= _GEN_7765;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_32 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_32 <= _GEN_2338;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_32 <= _GEN_7766;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_33 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_33 <= _GEN_2339;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_33 <= _GEN_7767;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_34 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_34 <= _GEN_2340;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_34 <= _GEN_7768;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_35 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_35 <= _GEN_2341;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_35 <= _GEN_7769;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_36 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_36 <= _GEN_2342;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_36 <= _GEN_7770;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_37 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_37 <= _GEN_2343;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_37 <= _GEN_7771;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_38 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_38 <= _GEN_2344;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_38 <= _GEN_7772;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_39 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_39 <= _GEN_2345;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_39 <= _GEN_7773;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_40 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_40 <= _GEN_2346;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_40 <= _GEN_7774;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_41 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_41 <= _GEN_2347;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_41 <= _GEN_7775;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_42 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_42 <= _GEN_2348;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_42 <= _GEN_7776;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_43 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_43 <= _GEN_2349;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_43 <= _GEN_7777;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_44 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_44 <= _GEN_2350;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_44 <= _GEN_7778;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_45 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_45 <= _GEN_2351;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_45 <= _GEN_7779;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_46 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_46 <= _GEN_2352;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_46 <= _GEN_7780;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_47 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_47 <= _GEN_2353;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_47 <= _GEN_7781;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_48 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_48 <= _GEN_2354;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_48 <= _GEN_7782;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_49 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_49 <= _GEN_2355;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_49 <= _GEN_7783;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_50 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_50 <= _GEN_2356;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_50 <= _GEN_7784;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_51 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_51 <= _GEN_2357;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_51 <= _GEN_7785;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_52 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_52 <= _GEN_2358;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_52 <= _GEN_7786;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_53 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_53 <= _GEN_2359;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_53 <= _GEN_7787;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_54 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_54 <= _GEN_2360;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_54 <= _GEN_7788;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_55 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_55 <= _GEN_2361;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_55 <= _GEN_7789;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_56 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_56 <= _GEN_2362;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_56 <= _GEN_7790;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_57 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_57 <= _GEN_2363;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_57 <= _GEN_7791;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_58 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_58 <= _GEN_2364;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_58 <= _GEN_7792;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_59 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_59 <= _GEN_2365;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_59 <= _GEN_7793;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_60 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_60 <= _GEN_2366;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_60 <= _GEN_7794;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_61 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_61 <= _GEN_2367;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_61 <= _GEN_7795;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_62 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_62 <= _GEN_2368;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_62 <= _GEN_7796;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_63 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_63 <= _GEN_2369;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_63 <= _GEN_7797;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_64 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_64 <= _GEN_2370;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_64 <= _GEN_7798;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_65 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_65 <= _GEN_2371;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_65 <= _GEN_7799;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_66 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_66 <= _GEN_2372;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_66 <= _GEN_7800;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_67 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_67 <= _GEN_2373;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_67 <= _GEN_7801;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_68 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_68 <= _GEN_2374;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_68 <= _GEN_7802;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_69 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_69 <= _GEN_2375;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_69 <= _GEN_7803;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_70 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_70 <= _GEN_2376;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_70 <= _GEN_7804;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_71 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_71 <= _GEN_2377;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_71 <= _GEN_7805;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_72 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_72 <= _GEN_2378;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_72 <= _GEN_7806;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_73 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_73 <= _GEN_2379;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_73 <= _GEN_7807;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_74 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_74 <= _GEN_2380;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_74 <= _GEN_7808;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_75 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_75 <= _GEN_2381;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_75 <= _GEN_7809;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_76 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_76 <= _GEN_2382;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_76 <= _GEN_7810;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_77 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_77 <= _GEN_2383;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_77 <= _GEN_7811;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_78 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_78 <= _GEN_2384;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_78 <= _GEN_7812;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_79 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_79 <= _GEN_2385;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_79 <= _GEN_7813;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_80 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_80 <= _GEN_2386;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_80 <= _GEN_7814;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_81 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_81 <= _GEN_2387;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_81 <= _GEN_7815;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_82 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_82 <= _GEN_2388;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_82 <= _GEN_7816;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_83 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_83 <= _GEN_2389;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_83 <= _GEN_7817;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_84 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_84 <= _GEN_2390;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_84 <= _GEN_7818;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_85 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_85 <= _GEN_2391;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_85 <= _GEN_7819;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_86 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_86 <= _GEN_2392;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_86 <= _GEN_7820;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_87 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_87 <= _GEN_2393;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_87 <= _GEN_7821;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_88 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_88 <= _GEN_2394;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_88 <= _GEN_7822;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_89 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_89 <= _GEN_2395;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_89 <= _GEN_7823;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_90 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_90 <= _GEN_2396;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_90 <= _GEN_7824;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_91 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_91 <= _GEN_2397;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_91 <= _GEN_7825;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_92 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_92 <= _GEN_2398;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_92 <= _GEN_7826;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_93 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_93 <= _GEN_2399;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_93 <= _GEN_7827;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_94 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_94 <= _GEN_2400;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_94 <= _GEN_7828;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_95 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_95 <= _GEN_2401;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_95 <= _GEN_7829;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_96 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_96 <= _GEN_2402;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_96 <= _GEN_7830;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_97 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_97 <= _GEN_2403;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_97 <= _GEN_7831;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_98 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_98 <= _GEN_2404;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_98 <= _GEN_7832;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_99 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_99 <= _GEN_2405;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_99 <= _GEN_7833;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_100 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_100 <= _GEN_2406;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_100 <= _GEN_7834;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_101 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_101 <= _GEN_2407;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_101 <= _GEN_7835;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_102 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_102 <= _GEN_2408;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_102 <= _GEN_7836;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_103 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_103 <= _GEN_2409;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_103 <= _GEN_7837;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_104 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_104 <= _GEN_2410;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_104 <= _GEN_7838;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_105 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_105 <= _GEN_2411;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_105 <= _GEN_7839;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_106 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_106 <= _GEN_2412;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_106 <= _GEN_7840;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_107 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_107 <= _GEN_2413;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_107 <= _GEN_7841;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_108 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_108 <= _GEN_2414;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_108 <= _GEN_7842;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_109 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_109 <= _GEN_2415;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_109 <= _GEN_7843;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_110 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_110 <= _GEN_2416;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_110 <= _GEN_7844;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_111 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_111 <= _GEN_2417;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_111 <= _GEN_7845;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_112 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_112 <= _GEN_2418;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_112 <= _GEN_7846;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_113 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_113 <= _GEN_2419;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_113 <= _GEN_7847;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_114 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_114 <= _GEN_2420;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_114 <= _GEN_7848;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_115 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_115 <= _GEN_2421;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_115 <= _GEN_7849;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_116 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_116 <= _GEN_2422;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_116 <= _GEN_7850;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_117 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_117 <= _GEN_2423;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_117 <= _GEN_7851;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_118 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_118 <= _GEN_2424;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_118 <= _GEN_7852;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_119 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_119 <= _GEN_2425;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_119 <= _GEN_7853;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_120 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_120 <= _GEN_2426;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_120 <= _GEN_7854;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_121 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_121 <= _GEN_2427;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_121 <= _GEN_7855;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_122 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_122 <= _GEN_2428;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_122 <= _GEN_7856;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_123 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_123 <= _GEN_2429;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_123 <= _GEN_7857;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_124 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_124 <= _GEN_2430;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_124 <= _GEN_7858;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_125 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_125 <= _GEN_2431;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_125 <= _GEN_7859;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_126 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_126 <= _GEN_2432;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_126 <= _GEN_7860;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_127 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_127 <= _GEN_2433;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_127 <= _GEN_7861;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_128 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_128 <= _GEN_2434;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_128 <= _GEN_7862;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_129 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_129 <= _GEN_2435;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_129 <= _GEN_7863;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_130 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_130 <= _GEN_2436;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_130 <= _GEN_7864;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_131 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_131 <= _GEN_2437;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_131 <= _GEN_7865;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_132 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_132 <= _GEN_2438;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_132 <= _GEN_7866;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_133 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_133 <= _GEN_2439;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_133 <= _GEN_7867;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_134 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_134 <= _GEN_2440;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_134 <= _GEN_7868;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_135 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_135 <= _GEN_2441;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_135 <= _GEN_7869;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_136 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_136 <= _GEN_2442;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_136 <= _GEN_7870;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_137 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_137 <= _GEN_2443;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_137 <= _GEN_7871;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_138 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_138 <= _GEN_2444;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_138 <= _GEN_7872;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_139 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_139 <= _GEN_2445;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_139 <= _GEN_7873;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_140 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_140 <= _GEN_2446;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_140 <= _GEN_7874;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_141 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_141 <= _GEN_2447;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_141 <= _GEN_7875;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_142 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_142 <= _GEN_2448;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_142 <= _GEN_7876;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_143 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_143 <= _GEN_2449;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_143 <= _GEN_7877;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_144 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_144 <= _GEN_2450;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_144 <= _GEN_7878;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_145 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_145 <= _GEN_2451;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_145 <= _GEN_7879;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_146 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_146 <= _GEN_2452;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_146 <= _GEN_7880;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_147 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_147 <= _GEN_2453;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_147 <= _GEN_7881;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_148 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_148 <= _GEN_2454;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_148 <= _GEN_7882;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_149 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_149 <= _GEN_2455;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_149 <= _GEN_7883;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_150 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_150 <= _GEN_2456;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_150 <= _GEN_7884;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_151 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_151 <= _GEN_2457;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_151 <= _GEN_7885;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_152 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_152 <= _GEN_2458;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_152 <= _GEN_7886;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_153 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_153 <= _GEN_2459;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_153 <= _GEN_7887;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_154 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_154 <= _GEN_2460;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_154 <= _GEN_7888;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_155 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_155 <= _GEN_2461;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_155 <= _GEN_7889;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_156 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_156 <= _GEN_2462;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_156 <= _GEN_7890;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_157 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_157 <= _GEN_2463;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_157 <= _GEN_7891;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_158 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_158 <= _GEN_2464;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_158 <= _GEN_7892;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_159 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_159 <= _GEN_2465;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_159 <= _GEN_7893;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_160 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_160 <= _GEN_2466;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_160 <= _GEN_7894;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_161 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_161 <= _GEN_2467;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_161 <= _GEN_7895;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_162 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_162 <= _GEN_2468;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_162 <= _GEN_7896;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_163 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_163 <= _GEN_2469;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_163 <= _GEN_7897;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_164 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_164 <= _GEN_2470;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_164 <= _GEN_7898;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_165 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_165 <= _GEN_2471;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_165 <= _GEN_7899;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_166 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_166 <= _GEN_2472;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_166 <= _GEN_7900;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_167 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_167 <= _GEN_2473;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_167 <= _GEN_7901;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_168 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_168 <= _GEN_2474;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_168 <= _GEN_7902;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_169 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_169 <= _GEN_2475;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_169 <= _GEN_7903;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_170 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_170 <= _GEN_2476;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_170 <= _GEN_7904;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_171 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_171 <= _GEN_2477;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_171 <= _GEN_7905;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_172 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_172 <= _GEN_2478;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_172 <= _GEN_7906;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_173 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_173 <= _GEN_2479;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_173 <= _GEN_7907;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_174 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_174 <= _GEN_2480;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_174 <= _GEN_7908;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_175 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_175 <= _GEN_2481;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_175 <= _GEN_7909;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_176 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_176 <= _GEN_2482;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_176 <= _GEN_7910;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_177 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_177 <= _GEN_2483;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_177 <= _GEN_7911;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_178 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_178 <= _GEN_2484;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_178 <= _GEN_7912;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_179 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_179 <= _GEN_2485;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_179 <= _GEN_7913;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_180 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_180 <= _GEN_2486;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_180 <= _GEN_7914;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_181 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_181 <= _GEN_2487;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_181 <= _GEN_7915;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_182 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_182 <= _GEN_2488;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_182 <= _GEN_7916;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_183 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_183 <= _GEN_2489;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_183 <= _GEN_7917;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_184 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_184 <= _GEN_2490;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_184 <= _GEN_7918;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_185 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_185 <= _GEN_2491;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_185 <= _GEN_7919;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_186 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_186 <= _GEN_2492;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_186 <= _GEN_7920;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_187 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_187 <= _GEN_2493;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_187 <= _GEN_7921;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_188 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_188 <= _GEN_2494;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_188 <= _GEN_7922;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_189 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_189 <= _GEN_2495;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_189 <= _GEN_7923;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_190 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_190 <= _GEN_2496;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_190 <= _GEN_7924;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_191 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_191 <= _GEN_2497;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_191 <= _GEN_7925;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_192 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_192 <= _GEN_2498;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_192 <= _GEN_7926;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_193 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_193 <= _GEN_2499;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_193 <= _GEN_7927;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_194 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_194 <= _GEN_2500;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_194 <= _GEN_7928;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_195 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_195 <= _GEN_2501;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_195 <= _GEN_7929;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_196 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_196 <= _GEN_2502;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_196 <= _GEN_7930;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_197 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_197 <= _GEN_2503;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_197 <= _GEN_7931;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_198 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_198 <= _GEN_2504;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_198 <= _GEN_7932;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_199 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_199 <= _GEN_2505;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_199 <= _GEN_7933;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_200 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_200 <= _GEN_2506;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_200 <= _GEN_7934;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_201 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_201 <= _GEN_2507;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_201 <= _GEN_7935;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_202 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_202 <= _GEN_2508;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_202 <= _GEN_7936;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_203 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_203 <= _GEN_2509;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_203 <= _GEN_7937;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_204 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_204 <= _GEN_2510;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_204 <= _GEN_7938;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_205 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_205 <= _GEN_2511;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_205 <= _GEN_7939;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_206 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_206 <= _GEN_2512;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_206 <= _GEN_7940;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_207 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_207 <= _GEN_2513;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_207 <= _GEN_7941;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_208 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_208 <= _GEN_2514;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_208 <= _GEN_7942;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_209 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_209 <= _GEN_2515;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_209 <= _GEN_7943;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_210 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_210 <= _GEN_2516;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_210 <= _GEN_7944;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_211 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_211 <= _GEN_2517;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_211 <= _GEN_7945;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_212 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_212 <= _GEN_2518;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_212 <= _GEN_7946;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_213 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_213 <= _GEN_2519;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_213 <= _GEN_7947;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_214 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_214 <= _GEN_2520;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_214 <= _GEN_7948;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_215 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_215 <= _GEN_2521;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_215 <= _GEN_7949;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_216 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_216 <= _GEN_2522;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_216 <= _GEN_7950;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_217 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_217 <= _GEN_2523;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_217 <= _GEN_7951;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_218 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_218 <= _GEN_2524;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_218 <= _GEN_7952;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_219 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_219 <= _GEN_2525;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_219 <= _GEN_7953;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_220 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_220 <= _GEN_2526;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_220 <= _GEN_7954;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_221 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_221 <= _GEN_2527;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_221 <= _GEN_7955;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_222 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_222 <= _GEN_2528;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_222 <= _GEN_7956;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_223 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_223 <= _GEN_2529;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_223 <= _GEN_7957;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_224 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_224 <= _GEN_2530;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_224 <= _GEN_7958;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_225 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_225 <= _GEN_2531;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_225 <= _GEN_7959;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_226 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_226 <= _GEN_2532;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_226 <= _GEN_7960;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_227 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_227 <= _GEN_2533;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_227 <= _GEN_7961;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_228 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_228 <= _GEN_2534;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_228 <= _GEN_7962;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_229 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_229 <= _GEN_2535;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_229 <= _GEN_7963;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_230 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_230 <= _GEN_2536;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_230 <= _GEN_7964;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_231 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_231 <= _GEN_2537;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_231 <= _GEN_7965;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_232 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_232 <= _GEN_2538;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_232 <= _GEN_7966;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_233 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_233 <= _GEN_2539;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_233 <= _GEN_7967;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_234 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_234 <= _GEN_2540;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_234 <= _GEN_7968;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_235 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_235 <= _GEN_2541;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_235 <= _GEN_7969;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_236 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_236 <= _GEN_2542;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_236 <= _GEN_7970;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_237 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_237 <= _GEN_2543;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_237 <= _GEN_7971;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_238 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_238 <= _GEN_2544;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_238 <= _GEN_7972;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_239 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_239 <= _GEN_2545;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_239 <= _GEN_7973;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_240 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_240 <= _GEN_2546;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_240 <= _GEN_7974;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_241 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_241 <= _GEN_2547;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_241 <= _GEN_7975;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_242 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_242 <= _GEN_2548;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_242 <= _GEN_7976;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_243 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_243 <= _GEN_2549;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_243 <= _GEN_7977;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_244 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_244 <= _GEN_2550;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_244 <= _GEN_7978;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_245 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_245 <= _GEN_2551;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_245 <= _GEN_7979;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_246 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_246 <= _GEN_2552;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_246 <= _GEN_7980;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_247 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_247 <= _GEN_2553;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_247 <= _GEN_7981;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_248 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_248 <= _GEN_2554;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_248 <= _GEN_7982;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_249 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_249 <= _GEN_2555;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_249 <= _GEN_7983;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_250 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_250 <= _GEN_2556;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_250 <= _GEN_7984;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_251 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_251 <= _GEN_2557;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_251 <= _GEN_7985;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_252 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_252 <= _GEN_2558;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_252 <= _GEN_7986;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_253 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_253 <= _GEN_2559;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_253 <= _GEN_7987;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_254 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_254 <= _GEN_2560;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_254 <= _GEN_7988;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_255 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          tag_255 <= _GEN_2561;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        tag_255 <= _GEN_7989;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_0 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_0 <= _GEN_2050;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_0 <= _GEN_7478;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_1 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_1 <= _GEN_2051;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_1 <= _GEN_7479;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_2 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_2 <= _GEN_2052;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_2 <= _GEN_7480;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_3 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_3 <= _GEN_2053;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_3 <= _GEN_7481;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_4 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_4 <= _GEN_2054;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_4 <= _GEN_7482;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_5 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_5 <= _GEN_2055;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_5 <= _GEN_7483;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_6 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_6 <= _GEN_2056;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_6 <= _GEN_7484;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_7 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_7 <= _GEN_2057;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_7 <= _GEN_7485;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_8 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_8 <= _GEN_2058;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_8 <= _GEN_7486;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_9 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_9 <= _GEN_2059;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_9 <= _GEN_7487;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_10 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_10 <= _GEN_2060;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_10 <= _GEN_7488;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_11 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_11 <= _GEN_2061;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_11 <= _GEN_7489;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_12 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_12 <= _GEN_2062;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_12 <= _GEN_7490;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_13 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_13 <= _GEN_2063;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_13 <= _GEN_7491;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_14 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_14 <= _GEN_2064;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_14 <= _GEN_7492;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_15 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_15 <= _GEN_2065;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_15 <= _GEN_7493;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_16 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_16 <= _GEN_2066;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_16 <= _GEN_7494;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_17 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_17 <= _GEN_2067;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_17 <= _GEN_7495;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_18 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_18 <= _GEN_2068;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_18 <= _GEN_7496;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_19 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_19 <= _GEN_2069;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_19 <= _GEN_7497;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_20 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_20 <= _GEN_2070;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_20 <= _GEN_7498;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_21 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_21 <= _GEN_2071;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_21 <= _GEN_7499;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_22 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_22 <= _GEN_2072;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_22 <= _GEN_7500;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_23 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_23 <= _GEN_2073;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_23 <= _GEN_7501;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_24 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_24 <= _GEN_2074;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_24 <= _GEN_7502;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_25 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_25 <= _GEN_2075;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_25 <= _GEN_7503;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_26 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_26 <= _GEN_2076;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_26 <= _GEN_7504;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_27 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_27 <= _GEN_2077;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_27 <= _GEN_7505;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_28 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_28 <= _GEN_2078;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_28 <= _GEN_7506;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_29 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_29 <= _GEN_2079;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_29 <= _GEN_7507;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_30 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_30 <= _GEN_2080;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_30 <= _GEN_7508;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_31 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_31 <= _GEN_2081;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_31 <= _GEN_7509;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_32 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_32 <= _GEN_2082;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_32 <= _GEN_7510;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_33 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_33 <= _GEN_2083;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_33 <= _GEN_7511;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_34 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_34 <= _GEN_2084;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_34 <= _GEN_7512;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_35 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_35 <= _GEN_2085;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_35 <= _GEN_7513;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_36 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_36 <= _GEN_2086;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_36 <= _GEN_7514;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_37 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_37 <= _GEN_2087;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_37 <= _GEN_7515;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_38 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_38 <= _GEN_2088;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_38 <= _GEN_7516;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_39 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_39 <= _GEN_2089;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_39 <= _GEN_7517;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_40 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_40 <= _GEN_2090;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_40 <= _GEN_7518;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_41 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_41 <= _GEN_2091;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_41 <= _GEN_7519;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_42 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_42 <= _GEN_2092;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_42 <= _GEN_7520;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_43 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_43 <= _GEN_2093;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_43 <= _GEN_7521;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_44 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_44 <= _GEN_2094;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_44 <= _GEN_7522;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_45 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_45 <= _GEN_2095;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_45 <= _GEN_7523;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_46 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_46 <= _GEN_2096;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_46 <= _GEN_7524;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_47 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_47 <= _GEN_2097;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_47 <= _GEN_7525;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_48 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_48 <= _GEN_2098;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_48 <= _GEN_7526;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_49 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_49 <= _GEN_2099;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_49 <= _GEN_7527;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_50 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_50 <= _GEN_2100;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_50 <= _GEN_7528;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_51 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_51 <= _GEN_2101;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_51 <= _GEN_7529;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_52 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_52 <= _GEN_2102;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_52 <= _GEN_7530;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_53 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_53 <= _GEN_2103;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_53 <= _GEN_7531;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_54 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_54 <= _GEN_2104;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_54 <= _GEN_7532;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_55 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_55 <= _GEN_2105;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_55 <= _GEN_7533;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_56 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_56 <= _GEN_2106;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_56 <= _GEN_7534;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_57 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_57 <= _GEN_2107;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_57 <= _GEN_7535;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_58 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_58 <= _GEN_2108;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_58 <= _GEN_7536;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_59 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_59 <= _GEN_2109;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_59 <= _GEN_7537;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_60 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_60 <= _GEN_2110;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_60 <= _GEN_7538;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_61 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_61 <= _GEN_2111;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_61 <= _GEN_7539;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_62 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_62 <= _GEN_2112;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_62 <= _GEN_7540;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_63 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_63 <= _GEN_2113;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_63 <= _GEN_7541;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_64 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_64 <= _GEN_2114;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_64 <= _GEN_7542;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_65 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_65 <= _GEN_2115;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_65 <= _GEN_7543;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_66 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_66 <= _GEN_2116;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_66 <= _GEN_7544;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_67 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_67 <= _GEN_2117;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_67 <= _GEN_7545;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_68 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_68 <= _GEN_2118;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_68 <= _GEN_7546;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_69 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_69 <= _GEN_2119;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_69 <= _GEN_7547;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_70 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_70 <= _GEN_2120;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_70 <= _GEN_7548;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_71 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_71 <= _GEN_2121;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_71 <= _GEN_7549;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_72 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_72 <= _GEN_2122;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_72 <= _GEN_7550;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_73 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_73 <= _GEN_2123;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_73 <= _GEN_7551;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_74 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_74 <= _GEN_2124;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_74 <= _GEN_7552;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_75 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_75 <= _GEN_2125;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_75 <= _GEN_7553;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_76 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_76 <= _GEN_2126;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_76 <= _GEN_7554;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_77 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_77 <= _GEN_2127;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_77 <= _GEN_7555;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_78 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_78 <= _GEN_2128;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_78 <= _GEN_7556;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_79 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_79 <= _GEN_2129;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_79 <= _GEN_7557;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_80 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_80 <= _GEN_2130;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_80 <= _GEN_7558;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_81 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_81 <= _GEN_2131;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_81 <= _GEN_7559;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_82 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_82 <= _GEN_2132;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_82 <= _GEN_7560;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_83 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_83 <= _GEN_2133;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_83 <= _GEN_7561;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_84 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_84 <= _GEN_2134;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_84 <= _GEN_7562;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_85 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_85 <= _GEN_2135;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_85 <= _GEN_7563;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_86 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_86 <= _GEN_2136;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_86 <= _GEN_7564;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_87 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_87 <= _GEN_2137;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_87 <= _GEN_7565;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_88 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_88 <= _GEN_2138;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_88 <= _GEN_7566;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_89 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_89 <= _GEN_2139;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_89 <= _GEN_7567;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_90 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_90 <= _GEN_2140;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_90 <= _GEN_7568;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_91 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_91 <= _GEN_2141;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_91 <= _GEN_7569;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_92 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_92 <= _GEN_2142;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_92 <= _GEN_7570;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_93 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_93 <= _GEN_2143;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_93 <= _GEN_7571;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_94 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_94 <= _GEN_2144;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_94 <= _GEN_7572;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_95 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_95 <= _GEN_2145;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_95 <= _GEN_7573;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_96 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_96 <= _GEN_2146;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_96 <= _GEN_7574;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_97 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_97 <= _GEN_2147;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_97 <= _GEN_7575;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_98 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_98 <= _GEN_2148;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_98 <= _GEN_7576;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_99 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_99 <= _GEN_2149;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_99 <= _GEN_7577;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_100 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_100 <= _GEN_2150;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_100 <= _GEN_7578;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_101 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_101 <= _GEN_2151;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_101 <= _GEN_7579;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_102 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_102 <= _GEN_2152;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_102 <= _GEN_7580;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_103 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_103 <= _GEN_2153;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_103 <= _GEN_7581;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_104 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_104 <= _GEN_2154;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_104 <= _GEN_7582;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_105 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_105 <= _GEN_2155;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_105 <= _GEN_7583;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_106 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_106 <= _GEN_2156;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_106 <= _GEN_7584;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_107 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_107 <= _GEN_2157;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_107 <= _GEN_7585;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_108 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_108 <= _GEN_2158;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_108 <= _GEN_7586;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_109 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_109 <= _GEN_2159;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_109 <= _GEN_7587;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_110 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_110 <= _GEN_2160;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_110 <= _GEN_7588;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_111 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_111 <= _GEN_2161;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_111 <= _GEN_7589;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_112 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_112 <= _GEN_2162;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_112 <= _GEN_7590;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_113 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_113 <= _GEN_2163;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_113 <= _GEN_7591;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_114 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_114 <= _GEN_2164;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_114 <= _GEN_7592;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_115 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_115 <= _GEN_2165;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_115 <= _GEN_7593;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_116 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_116 <= _GEN_2166;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_116 <= _GEN_7594;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_117 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_117 <= _GEN_2167;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_117 <= _GEN_7595;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_118 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_118 <= _GEN_2168;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_118 <= _GEN_7596;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_119 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_119 <= _GEN_2169;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_119 <= _GEN_7597;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_120 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_120 <= _GEN_2170;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_120 <= _GEN_7598;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_121 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_121 <= _GEN_2171;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_121 <= _GEN_7599;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_122 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_122 <= _GEN_2172;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_122 <= _GEN_7600;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_123 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_123 <= _GEN_2173;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_123 <= _GEN_7601;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_124 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_124 <= _GEN_2174;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_124 <= _GEN_7602;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_125 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_125 <= _GEN_2175;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_125 <= _GEN_7603;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_126 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_126 <= _GEN_2176;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_126 <= _GEN_7604;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_127 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_127 <= _GEN_2177;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_127 <= _GEN_7605;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_128 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_128 <= _GEN_2178;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_128 <= _GEN_7606;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_129 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_129 <= _GEN_2179;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_129 <= _GEN_7607;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_130 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_130 <= _GEN_2180;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_130 <= _GEN_7608;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_131 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_131 <= _GEN_2181;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_131 <= _GEN_7609;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_132 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_132 <= _GEN_2182;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_132 <= _GEN_7610;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_133 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_133 <= _GEN_2183;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_133 <= _GEN_7611;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_134 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_134 <= _GEN_2184;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_134 <= _GEN_7612;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_135 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_135 <= _GEN_2185;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_135 <= _GEN_7613;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_136 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_136 <= _GEN_2186;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_136 <= _GEN_7614;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_137 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_137 <= _GEN_2187;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_137 <= _GEN_7615;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_138 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_138 <= _GEN_2188;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_138 <= _GEN_7616;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_139 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_139 <= _GEN_2189;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_139 <= _GEN_7617;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_140 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_140 <= _GEN_2190;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_140 <= _GEN_7618;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_141 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_141 <= _GEN_2191;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_141 <= _GEN_7619;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_142 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_142 <= _GEN_2192;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_142 <= _GEN_7620;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_143 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_143 <= _GEN_2193;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_143 <= _GEN_7621;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_144 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_144 <= _GEN_2194;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_144 <= _GEN_7622;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_145 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_145 <= _GEN_2195;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_145 <= _GEN_7623;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_146 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_146 <= _GEN_2196;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_146 <= _GEN_7624;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_147 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_147 <= _GEN_2197;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_147 <= _GEN_7625;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_148 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_148 <= _GEN_2198;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_148 <= _GEN_7626;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_149 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_149 <= _GEN_2199;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_149 <= _GEN_7627;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_150 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_150 <= _GEN_2200;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_150 <= _GEN_7628;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_151 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_151 <= _GEN_2201;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_151 <= _GEN_7629;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_152 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_152 <= _GEN_2202;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_152 <= _GEN_7630;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_153 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_153 <= _GEN_2203;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_153 <= _GEN_7631;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_154 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_154 <= _GEN_2204;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_154 <= _GEN_7632;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_155 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_155 <= _GEN_2205;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_155 <= _GEN_7633;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_156 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_156 <= _GEN_2206;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_156 <= _GEN_7634;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_157 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_157 <= _GEN_2207;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_157 <= _GEN_7635;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_158 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_158 <= _GEN_2208;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_158 <= _GEN_7636;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_159 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_159 <= _GEN_2209;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_159 <= _GEN_7637;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_160 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_160 <= _GEN_2210;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_160 <= _GEN_7638;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_161 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_161 <= _GEN_2211;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_161 <= _GEN_7639;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_162 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_162 <= _GEN_2212;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_162 <= _GEN_7640;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_163 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_163 <= _GEN_2213;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_163 <= _GEN_7641;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_164 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_164 <= _GEN_2214;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_164 <= _GEN_7642;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_165 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_165 <= _GEN_2215;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_165 <= _GEN_7643;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_166 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_166 <= _GEN_2216;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_166 <= _GEN_7644;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_167 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_167 <= _GEN_2217;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_167 <= _GEN_7645;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_168 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_168 <= _GEN_2218;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_168 <= _GEN_7646;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_169 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_169 <= _GEN_2219;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_169 <= _GEN_7647;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_170 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_170 <= _GEN_2220;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_170 <= _GEN_7648;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_171 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_171 <= _GEN_2221;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_171 <= _GEN_7649;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_172 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_172 <= _GEN_2222;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_172 <= _GEN_7650;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_173 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_173 <= _GEN_2223;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_173 <= _GEN_7651;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_174 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_174 <= _GEN_2224;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_174 <= _GEN_7652;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_175 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_175 <= _GEN_2225;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_175 <= _GEN_7653;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_176 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_176 <= _GEN_2226;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_176 <= _GEN_7654;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_177 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_177 <= _GEN_2227;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_177 <= _GEN_7655;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_178 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_178 <= _GEN_2228;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_178 <= _GEN_7656;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_179 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_179 <= _GEN_2229;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_179 <= _GEN_7657;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_180 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_180 <= _GEN_2230;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_180 <= _GEN_7658;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_181 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_181 <= _GEN_2231;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_181 <= _GEN_7659;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_182 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_182 <= _GEN_2232;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_182 <= _GEN_7660;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_183 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_183 <= _GEN_2233;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_183 <= _GEN_7661;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_184 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_184 <= _GEN_2234;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_184 <= _GEN_7662;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_185 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_185 <= _GEN_2235;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_185 <= _GEN_7663;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_186 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_186 <= _GEN_2236;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_186 <= _GEN_7664;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_187 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_187 <= _GEN_2237;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_187 <= _GEN_7665;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_188 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_188 <= _GEN_2238;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_188 <= _GEN_7666;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_189 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_189 <= _GEN_2239;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_189 <= _GEN_7667;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_190 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_190 <= _GEN_2240;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_190 <= _GEN_7668;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_191 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_191 <= _GEN_2241;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_191 <= _GEN_7669;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_192 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_192 <= _GEN_2242;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_192 <= _GEN_7670;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_193 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_193 <= _GEN_2243;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_193 <= _GEN_7671;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_194 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_194 <= _GEN_2244;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_194 <= _GEN_7672;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_195 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_195 <= _GEN_2245;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_195 <= _GEN_7673;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_196 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_196 <= _GEN_2246;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_196 <= _GEN_7674;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_197 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_197 <= _GEN_2247;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_197 <= _GEN_7675;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_198 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_198 <= _GEN_2248;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_198 <= _GEN_7676;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_199 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_199 <= _GEN_2249;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_199 <= _GEN_7677;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_200 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_200 <= _GEN_2250;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_200 <= _GEN_7678;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_201 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_201 <= _GEN_2251;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_201 <= _GEN_7679;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_202 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_202 <= _GEN_2252;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_202 <= _GEN_7680;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_203 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_203 <= _GEN_2253;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_203 <= _GEN_7681;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_204 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_204 <= _GEN_2254;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_204 <= _GEN_7682;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_205 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_205 <= _GEN_2255;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_205 <= _GEN_7683;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_206 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_206 <= _GEN_2256;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_206 <= _GEN_7684;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_207 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_207 <= _GEN_2257;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_207 <= _GEN_7685;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_208 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_208 <= _GEN_2258;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_208 <= _GEN_7686;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_209 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_209 <= _GEN_2259;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_209 <= _GEN_7687;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_210 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_210 <= _GEN_2260;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_210 <= _GEN_7688;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_211 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_211 <= _GEN_2261;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_211 <= _GEN_7689;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_212 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_212 <= _GEN_2262;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_212 <= _GEN_7690;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_213 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_213 <= _GEN_2263;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_213 <= _GEN_7691;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_214 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_214 <= _GEN_2264;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_214 <= _GEN_7692;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_215 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_215 <= _GEN_2265;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_215 <= _GEN_7693;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_216 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_216 <= _GEN_2266;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_216 <= _GEN_7694;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_217 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_217 <= _GEN_2267;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_217 <= _GEN_7695;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_218 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_218 <= _GEN_2268;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_218 <= _GEN_7696;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_219 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_219 <= _GEN_2269;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_219 <= _GEN_7697;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_220 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_220 <= _GEN_2270;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_220 <= _GEN_7698;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_221 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_221 <= _GEN_2271;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_221 <= _GEN_7699;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_222 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_222 <= _GEN_2272;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_222 <= _GEN_7700;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_223 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_223 <= _GEN_2273;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_223 <= _GEN_7701;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_224 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_224 <= _GEN_2274;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_224 <= _GEN_7702;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_225 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_225 <= _GEN_2275;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_225 <= _GEN_7703;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_226 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_226 <= _GEN_2276;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_226 <= _GEN_7704;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_227 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_227 <= _GEN_2277;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_227 <= _GEN_7705;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_228 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_228 <= _GEN_2278;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_228 <= _GEN_7706;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_229 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_229 <= _GEN_2279;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_229 <= _GEN_7707;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_230 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_230 <= _GEN_2280;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_230 <= _GEN_7708;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_231 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_231 <= _GEN_2281;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_231 <= _GEN_7709;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_232 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_232 <= _GEN_2282;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_232 <= _GEN_7710;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_233 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_233 <= _GEN_2283;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_233 <= _GEN_7711;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_234 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_234 <= _GEN_2284;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_234 <= _GEN_7712;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_235 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_235 <= _GEN_2285;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_235 <= _GEN_7713;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_236 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_236 <= _GEN_2286;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_236 <= _GEN_7714;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_237 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_237 <= _GEN_2287;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_237 <= _GEN_7715;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_238 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_238 <= _GEN_2288;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_238 <= _GEN_7716;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_239 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_239 <= _GEN_2289;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_239 <= _GEN_7717;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_240 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_240 <= _GEN_2290;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_240 <= _GEN_7718;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_241 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_241 <= _GEN_2291;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_241 <= _GEN_7719;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_242 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_242 <= _GEN_2292;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_242 <= _GEN_7720;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_243 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_243 <= _GEN_2293;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_243 <= _GEN_7721;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_244 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_244 <= _GEN_2294;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_244 <= _GEN_7722;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_245 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_245 <= _GEN_2295;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_245 <= _GEN_7723;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_246 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_246 <= _GEN_2296;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_246 <= _GEN_7724;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_247 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_247 <= _GEN_2297;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_247 <= _GEN_7725;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_248 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_248 <= _GEN_2298;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_248 <= _GEN_7726;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_249 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_249 <= _GEN_2299;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_249 <= _GEN_7727;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_250 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_250 <= _GEN_2300;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_250 <= _GEN_7728;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_251 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_251 <= _GEN_2301;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_251 <= _GEN_7729;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_252 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_252 <= _GEN_2302;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_252 <= _GEN_7730;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_253 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_253 <= _GEN_2303;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_253 <= _GEN_7731;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_254 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_254 <= _GEN_2304;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_254 <= _GEN_7732;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_255 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          valid_255 <= _GEN_2305;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        valid_255 <= _GEN_7733;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_0 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_0 <= _GEN_2822;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_0 <= _GEN_7990;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_1 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_1 <= _GEN_2823;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_1 <= _GEN_7991;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_2 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_2 <= _GEN_2824;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_2 <= _GEN_7992;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_3 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_3 <= _GEN_2825;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_3 <= _GEN_7993;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_4 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_4 <= _GEN_2826;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_4 <= _GEN_7994;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_5 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_5 <= _GEN_2827;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_5 <= _GEN_7995;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_6 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_6 <= _GEN_2828;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_6 <= _GEN_7996;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_7 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_7 <= _GEN_2829;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_7 <= _GEN_7997;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_8 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_8 <= _GEN_2830;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_8 <= _GEN_7998;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_9 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_9 <= _GEN_2831;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_9 <= _GEN_7999;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_10 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_10 <= _GEN_2832;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_10 <= _GEN_8000;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_11 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_11 <= _GEN_2833;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_11 <= _GEN_8001;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_12 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_12 <= _GEN_2834;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_12 <= _GEN_8002;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_13 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_13 <= _GEN_2835;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_13 <= _GEN_8003;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_14 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_14 <= _GEN_2836;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_14 <= _GEN_8004;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_15 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_15 <= _GEN_2837;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_15 <= _GEN_8005;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_16 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_16 <= _GEN_2838;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_16 <= _GEN_8006;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_17 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_17 <= _GEN_2839;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_17 <= _GEN_8007;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_18 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_18 <= _GEN_2840;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_18 <= _GEN_8008;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_19 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_19 <= _GEN_2841;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_19 <= _GEN_8009;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_20 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_20 <= _GEN_2842;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_20 <= _GEN_8010;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_21 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_21 <= _GEN_2843;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_21 <= _GEN_8011;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_22 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_22 <= _GEN_2844;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_22 <= _GEN_8012;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_23 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_23 <= _GEN_2845;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_23 <= _GEN_8013;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_24 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_24 <= _GEN_2846;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_24 <= _GEN_8014;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_25 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_25 <= _GEN_2847;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_25 <= _GEN_8015;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_26 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_26 <= _GEN_2848;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_26 <= _GEN_8016;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_27 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_27 <= _GEN_2849;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_27 <= _GEN_8017;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_28 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_28 <= _GEN_2850;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_28 <= _GEN_8018;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_29 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_29 <= _GEN_2851;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_29 <= _GEN_8019;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_30 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_30 <= _GEN_2852;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_30 <= _GEN_8020;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_31 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_31 <= _GEN_2853;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_31 <= _GEN_8021;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_32 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_32 <= _GEN_2854;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_32 <= _GEN_8022;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_33 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_33 <= _GEN_2855;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_33 <= _GEN_8023;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_34 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_34 <= _GEN_2856;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_34 <= _GEN_8024;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_35 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_35 <= _GEN_2857;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_35 <= _GEN_8025;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_36 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_36 <= _GEN_2858;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_36 <= _GEN_8026;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_37 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_37 <= _GEN_2859;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_37 <= _GEN_8027;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_38 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_38 <= _GEN_2860;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_38 <= _GEN_8028;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_39 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_39 <= _GEN_2861;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_39 <= _GEN_8029;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_40 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_40 <= _GEN_2862;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_40 <= _GEN_8030;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_41 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_41 <= _GEN_2863;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_41 <= _GEN_8031;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_42 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_42 <= _GEN_2864;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_42 <= _GEN_8032;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_43 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_43 <= _GEN_2865;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_43 <= _GEN_8033;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_44 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_44 <= _GEN_2866;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_44 <= _GEN_8034;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_45 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_45 <= _GEN_2867;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_45 <= _GEN_8035;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_46 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_46 <= _GEN_2868;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_46 <= _GEN_8036;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_47 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_47 <= _GEN_2869;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_47 <= _GEN_8037;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_48 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_48 <= _GEN_2870;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_48 <= _GEN_8038;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_49 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_49 <= _GEN_2871;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_49 <= _GEN_8039;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_50 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_50 <= _GEN_2872;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_50 <= _GEN_8040;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_51 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_51 <= _GEN_2873;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_51 <= _GEN_8041;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_52 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_52 <= _GEN_2874;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_52 <= _GEN_8042;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_53 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_53 <= _GEN_2875;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_53 <= _GEN_8043;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_54 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_54 <= _GEN_2876;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_54 <= _GEN_8044;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_55 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_55 <= _GEN_2877;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_55 <= _GEN_8045;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_56 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_56 <= _GEN_2878;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_56 <= _GEN_8046;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_57 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_57 <= _GEN_2879;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_57 <= _GEN_8047;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_58 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_58 <= _GEN_2880;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_58 <= _GEN_8048;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_59 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_59 <= _GEN_2881;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_59 <= _GEN_8049;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_60 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_60 <= _GEN_2882;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_60 <= _GEN_8050;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_61 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_61 <= _GEN_2883;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_61 <= _GEN_8051;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_62 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_62 <= _GEN_2884;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_62 <= _GEN_8052;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_63 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_63 <= _GEN_2885;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_63 <= _GEN_8053;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_64 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_64 <= _GEN_2886;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_64 <= _GEN_8054;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_65 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_65 <= _GEN_2887;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_65 <= _GEN_8055;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_66 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_66 <= _GEN_2888;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_66 <= _GEN_8056;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_67 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_67 <= _GEN_2889;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_67 <= _GEN_8057;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_68 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_68 <= _GEN_2890;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_68 <= _GEN_8058;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_69 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_69 <= _GEN_2891;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_69 <= _GEN_8059;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_70 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_70 <= _GEN_2892;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_70 <= _GEN_8060;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_71 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_71 <= _GEN_2893;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_71 <= _GEN_8061;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_72 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_72 <= _GEN_2894;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_72 <= _GEN_8062;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_73 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_73 <= _GEN_2895;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_73 <= _GEN_8063;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_74 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_74 <= _GEN_2896;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_74 <= _GEN_8064;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_75 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_75 <= _GEN_2897;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_75 <= _GEN_8065;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_76 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_76 <= _GEN_2898;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_76 <= _GEN_8066;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_77 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_77 <= _GEN_2899;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_77 <= _GEN_8067;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_78 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_78 <= _GEN_2900;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_78 <= _GEN_8068;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_79 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_79 <= _GEN_2901;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_79 <= _GEN_8069;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_80 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_80 <= _GEN_2902;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_80 <= _GEN_8070;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_81 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_81 <= _GEN_2903;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_81 <= _GEN_8071;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_82 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_82 <= _GEN_2904;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_82 <= _GEN_8072;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_83 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_83 <= _GEN_2905;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_83 <= _GEN_8073;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_84 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_84 <= _GEN_2906;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_84 <= _GEN_8074;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_85 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_85 <= _GEN_2907;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_85 <= _GEN_8075;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_86 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_86 <= _GEN_2908;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_86 <= _GEN_8076;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_87 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_87 <= _GEN_2909;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_87 <= _GEN_8077;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_88 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_88 <= _GEN_2910;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_88 <= _GEN_8078;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_89 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_89 <= _GEN_2911;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_89 <= _GEN_8079;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_90 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_90 <= _GEN_2912;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_90 <= _GEN_8080;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_91 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_91 <= _GEN_2913;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_91 <= _GEN_8081;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_92 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_92 <= _GEN_2914;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_92 <= _GEN_8082;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_93 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_93 <= _GEN_2915;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_93 <= _GEN_8083;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_94 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_94 <= _GEN_2916;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_94 <= _GEN_8084;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_95 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_95 <= _GEN_2917;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_95 <= _GEN_8085;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_96 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_96 <= _GEN_2918;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_96 <= _GEN_8086;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_97 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_97 <= _GEN_2919;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_97 <= _GEN_8087;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_98 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_98 <= _GEN_2920;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_98 <= _GEN_8088;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_99 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_99 <= _GEN_2921;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_99 <= _GEN_8089;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_100 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_100 <= _GEN_2922;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_100 <= _GEN_8090;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_101 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_101 <= _GEN_2923;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_101 <= _GEN_8091;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_102 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_102 <= _GEN_2924;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_102 <= _GEN_8092;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_103 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_103 <= _GEN_2925;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_103 <= _GEN_8093;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_104 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_104 <= _GEN_2926;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_104 <= _GEN_8094;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_105 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_105 <= _GEN_2927;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_105 <= _GEN_8095;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_106 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_106 <= _GEN_2928;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_106 <= _GEN_8096;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_107 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_107 <= _GEN_2929;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_107 <= _GEN_8097;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_108 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_108 <= _GEN_2930;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_108 <= _GEN_8098;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_109 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_109 <= _GEN_2931;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_109 <= _GEN_8099;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_110 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_110 <= _GEN_2932;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_110 <= _GEN_8100;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_111 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_111 <= _GEN_2933;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_111 <= _GEN_8101;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_112 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_112 <= _GEN_2934;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_112 <= _GEN_8102;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_113 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_113 <= _GEN_2935;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_113 <= _GEN_8103;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_114 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_114 <= _GEN_2936;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_114 <= _GEN_8104;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_115 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_115 <= _GEN_2937;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_115 <= _GEN_8105;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_116 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_116 <= _GEN_2938;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_116 <= _GEN_8106;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_117 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_117 <= _GEN_2939;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_117 <= _GEN_8107;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_118 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_118 <= _GEN_2940;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_118 <= _GEN_8108;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_119 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_119 <= _GEN_2941;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_119 <= _GEN_8109;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_120 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_120 <= _GEN_2942;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_120 <= _GEN_8110;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_121 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_121 <= _GEN_2943;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_121 <= _GEN_8111;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_122 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_122 <= _GEN_2944;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_122 <= _GEN_8112;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_123 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_123 <= _GEN_2945;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_123 <= _GEN_8113;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_124 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_124 <= _GEN_2946;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_124 <= _GEN_8114;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_125 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_125 <= _GEN_2947;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_125 <= _GEN_8115;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_126 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_126 <= _GEN_2948;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_126 <= _GEN_8116;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_127 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_127 <= _GEN_2949;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_127 <= _GEN_8117;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_128 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_128 <= _GEN_2950;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_128 <= _GEN_8118;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_129 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_129 <= _GEN_2951;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_129 <= _GEN_8119;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_130 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_130 <= _GEN_2952;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_130 <= _GEN_8120;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_131 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_131 <= _GEN_2953;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_131 <= _GEN_8121;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_132 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_132 <= _GEN_2954;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_132 <= _GEN_8122;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_133 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_133 <= _GEN_2955;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_133 <= _GEN_8123;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_134 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_134 <= _GEN_2956;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_134 <= _GEN_8124;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_135 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_135 <= _GEN_2957;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_135 <= _GEN_8125;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_136 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_136 <= _GEN_2958;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_136 <= _GEN_8126;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_137 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_137 <= _GEN_2959;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_137 <= _GEN_8127;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_138 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_138 <= _GEN_2960;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_138 <= _GEN_8128;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_139 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_139 <= _GEN_2961;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_139 <= _GEN_8129;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_140 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_140 <= _GEN_2962;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_140 <= _GEN_8130;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_141 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_141 <= _GEN_2963;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_141 <= _GEN_8131;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_142 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_142 <= _GEN_2964;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_142 <= _GEN_8132;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_143 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_143 <= _GEN_2965;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_143 <= _GEN_8133;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_144 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_144 <= _GEN_2966;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_144 <= _GEN_8134;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_145 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_145 <= _GEN_2967;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_145 <= _GEN_8135;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_146 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_146 <= _GEN_2968;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_146 <= _GEN_8136;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_147 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_147 <= _GEN_2969;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_147 <= _GEN_8137;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_148 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_148 <= _GEN_2970;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_148 <= _GEN_8138;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_149 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_149 <= _GEN_2971;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_149 <= _GEN_8139;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_150 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_150 <= _GEN_2972;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_150 <= _GEN_8140;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_151 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_151 <= _GEN_2973;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_151 <= _GEN_8141;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_152 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_152 <= _GEN_2974;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_152 <= _GEN_8142;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_153 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_153 <= _GEN_2975;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_153 <= _GEN_8143;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_154 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_154 <= _GEN_2976;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_154 <= _GEN_8144;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_155 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_155 <= _GEN_2977;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_155 <= _GEN_8145;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_156 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_156 <= _GEN_2978;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_156 <= _GEN_8146;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_157 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_157 <= _GEN_2979;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_157 <= _GEN_8147;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_158 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_158 <= _GEN_2980;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_158 <= _GEN_8148;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_159 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_159 <= _GEN_2981;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_159 <= _GEN_8149;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_160 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_160 <= _GEN_2982;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_160 <= _GEN_8150;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_161 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_161 <= _GEN_2983;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_161 <= _GEN_8151;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_162 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_162 <= _GEN_2984;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_162 <= _GEN_8152;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_163 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_163 <= _GEN_2985;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_163 <= _GEN_8153;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_164 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_164 <= _GEN_2986;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_164 <= _GEN_8154;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_165 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_165 <= _GEN_2987;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_165 <= _GEN_8155;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_166 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_166 <= _GEN_2988;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_166 <= _GEN_8156;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_167 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_167 <= _GEN_2989;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_167 <= _GEN_8157;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_168 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_168 <= _GEN_2990;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_168 <= _GEN_8158;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_169 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_169 <= _GEN_2991;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_169 <= _GEN_8159;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_170 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_170 <= _GEN_2992;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_170 <= _GEN_8160;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_171 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_171 <= _GEN_2993;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_171 <= _GEN_8161;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_172 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_172 <= _GEN_2994;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_172 <= _GEN_8162;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_173 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_173 <= _GEN_2995;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_173 <= _GEN_8163;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_174 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_174 <= _GEN_2996;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_174 <= _GEN_8164;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_175 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_175 <= _GEN_2997;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_175 <= _GEN_8165;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_176 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_176 <= _GEN_2998;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_176 <= _GEN_8166;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_177 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_177 <= _GEN_2999;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_177 <= _GEN_8167;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_178 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_178 <= _GEN_3000;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_178 <= _GEN_8168;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_179 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_179 <= _GEN_3001;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_179 <= _GEN_8169;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_180 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_180 <= _GEN_3002;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_180 <= _GEN_8170;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_181 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_181 <= _GEN_3003;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_181 <= _GEN_8171;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_182 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_182 <= _GEN_3004;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_182 <= _GEN_8172;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_183 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_183 <= _GEN_3005;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_183 <= _GEN_8173;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_184 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_184 <= _GEN_3006;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_184 <= _GEN_8174;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_185 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_185 <= _GEN_3007;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_185 <= _GEN_8175;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_186 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_186 <= _GEN_3008;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_186 <= _GEN_8176;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_187 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_187 <= _GEN_3009;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_187 <= _GEN_8177;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_188 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_188 <= _GEN_3010;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_188 <= _GEN_8178;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_189 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_189 <= _GEN_3011;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_189 <= _GEN_8179;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_190 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_190 <= _GEN_3012;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_190 <= _GEN_8180;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_191 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_191 <= _GEN_3013;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_191 <= _GEN_8181;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_192 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_192 <= _GEN_3014;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_192 <= _GEN_8182;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_193 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_193 <= _GEN_3015;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_193 <= _GEN_8183;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_194 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_194 <= _GEN_3016;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_194 <= _GEN_8184;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_195 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_195 <= _GEN_3017;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_195 <= _GEN_8185;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_196 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_196 <= _GEN_3018;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_196 <= _GEN_8186;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_197 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_197 <= _GEN_3019;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_197 <= _GEN_8187;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_198 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_198 <= _GEN_3020;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_198 <= _GEN_8188;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_199 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_199 <= _GEN_3021;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_199 <= _GEN_8189;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_200 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_200 <= _GEN_3022;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_200 <= _GEN_8190;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_201 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_201 <= _GEN_3023;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_201 <= _GEN_8191;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_202 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_202 <= _GEN_3024;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_202 <= _GEN_8192;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_203 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_203 <= _GEN_3025;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_203 <= _GEN_8193;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_204 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_204 <= _GEN_3026;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_204 <= _GEN_8194;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_205 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_205 <= _GEN_3027;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_205 <= _GEN_8195;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_206 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_206 <= _GEN_3028;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_206 <= _GEN_8196;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_207 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_207 <= _GEN_3029;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_207 <= _GEN_8197;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_208 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_208 <= _GEN_3030;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_208 <= _GEN_8198;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_209 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_209 <= _GEN_3031;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_209 <= _GEN_8199;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_210 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_210 <= _GEN_3032;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_210 <= _GEN_8200;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_211 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_211 <= _GEN_3033;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_211 <= _GEN_8201;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_212 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_212 <= _GEN_3034;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_212 <= _GEN_8202;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_213 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_213 <= _GEN_3035;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_213 <= _GEN_8203;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_214 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_214 <= _GEN_3036;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_214 <= _GEN_8204;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_215 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_215 <= _GEN_3037;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_215 <= _GEN_8205;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_216 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_216 <= _GEN_3038;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_216 <= _GEN_8206;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_217 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_217 <= _GEN_3039;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_217 <= _GEN_8207;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_218 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_218 <= _GEN_3040;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_218 <= _GEN_8208;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_219 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_219 <= _GEN_3041;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_219 <= _GEN_8209;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_220 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_220 <= _GEN_3042;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_220 <= _GEN_8210;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_221 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_221 <= _GEN_3043;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_221 <= _GEN_8211;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_222 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_222 <= _GEN_3044;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_222 <= _GEN_8212;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_223 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_223 <= _GEN_3045;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_223 <= _GEN_8213;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_224 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_224 <= _GEN_3046;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_224 <= _GEN_8214;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_225 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_225 <= _GEN_3047;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_225 <= _GEN_8215;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_226 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_226 <= _GEN_3048;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_226 <= _GEN_8216;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_227 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_227 <= _GEN_3049;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_227 <= _GEN_8217;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_228 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_228 <= _GEN_3050;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_228 <= _GEN_8218;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_229 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_229 <= _GEN_3051;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_229 <= _GEN_8219;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_230 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_230 <= _GEN_3052;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_230 <= _GEN_8220;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_231 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_231 <= _GEN_3053;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_231 <= _GEN_8221;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_232 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_232 <= _GEN_3054;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_232 <= _GEN_8222;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_233 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_233 <= _GEN_3055;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_233 <= _GEN_8223;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_234 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_234 <= _GEN_3056;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_234 <= _GEN_8224;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_235 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_235 <= _GEN_3057;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_235 <= _GEN_8225;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_236 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_236 <= _GEN_3058;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_236 <= _GEN_8226;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_237 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_237 <= _GEN_3059;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_237 <= _GEN_8227;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_238 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_238 <= _GEN_3060;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_238 <= _GEN_8228;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_239 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_239 <= _GEN_3061;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_239 <= _GEN_8229;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_240 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_240 <= _GEN_3062;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_240 <= _GEN_8230;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_241 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_241 <= _GEN_3063;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_241 <= _GEN_8231;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_242 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_242 <= _GEN_3064;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_242 <= _GEN_8232;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_243 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_243 <= _GEN_3065;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_243 <= _GEN_8233;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_244 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_244 <= _GEN_3066;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_244 <= _GEN_8234;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_245 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_245 <= _GEN_3067;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_245 <= _GEN_8235;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_246 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_246 <= _GEN_3068;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_246 <= _GEN_8236;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_247 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_247 <= _GEN_3069;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_247 <= _GEN_8237;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_248 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_248 <= _GEN_3070;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_248 <= _GEN_8238;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_249 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_249 <= _GEN_3071;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_249 <= _GEN_8239;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_250 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_250 <= _GEN_3072;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_250 <= _GEN_8240;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_251 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_251 <= _GEN_3073;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_251 <= _GEN_8241;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_252 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_252 <= _GEN_3074;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_252 <= _GEN_8242;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_253 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_253 <= _GEN_3075;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_253 <= _GEN_8243;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_254 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_254 <= _GEN_3076;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_254 <= _GEN_8244;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_255 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          dirty_255 <= _GEN_3077;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        dirty_255 <= _GEN_8245;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_0 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_0 <= _GEN_2562;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_0 <= _GEN_8246;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_1 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_1 <= _GEN_2563;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_1 <= _GEN_8247;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_2 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_2 <= _GEN_2564;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_2 <= _GEN_8248;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_3 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_3 <= _GEN_2565;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_3 <= _GEN_8249;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_4 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_4 <= _GEN_2566;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_4 <= _GEN_8250;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_5 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_5 <= _GEN_2567;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_5 <= _GEN_8251;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_6 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_6 <= _GEN_2568;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_6 <= _GEN_8252;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_7 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_7 <= _GEN_2569;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_7 <= _GEN_8253;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_8 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_8 <= _GEN_2570;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_8 <= _GEN_8254;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_9 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_9 <= _GEN_2571;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_9 <= _GEN_8255;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_10 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_10 <= _GEN_2572;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_10 <= _GEN_8256;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_11 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_11 <= _GEN_2573;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_11 <= _GEN_8257;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_12 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_12 <= _GEN_2574;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_12 <= _GEN_8258;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_13 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_13 <= _GEN_2575;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_13 <= _GEN_8259;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_14 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_14 <= _GEN_2576;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_14 <= _GEN_8260;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_15 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_15 <= _GEN_2577;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_15 <= _GEN_8261;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_16 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_16 <= _GEN_2578;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_16 <= _GEN_8262;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_17 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_17 <= _GEN_2579;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_17 <= _GEN_8263;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_18 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_18 <= _GEN_2580;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_18 <= _GEN_8264;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_19 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_19 <= _GEN_2581;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_19 <= _GEN_8265;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_20 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_20 <= _GEN_2582;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_20 <= _GEN_8266;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_21 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_21 <= _GEN_2583;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_21 <= _GEN_8267;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_22 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_22 <= _GEN_2584;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_22 <= _GEN_8268;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_23 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_23 <= _GEN_2585;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_23 <= _GEN_8269;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_24 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_24 <= _GEN_2586;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_24 <= _GEN_8270;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_25 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_25 <= _GEN_2587;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_25 <= _GEN_8271;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_26 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_26 <= _GEN_2588;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_26 <= _GEN_8272;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_27 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_27 <= _GEN_2589;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_27 <= _GEN_8273;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_28 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_28 <= _GEN_2590;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_28 <= _GEN_8274;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_29 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_29 <= _GEN_2591;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_29 <= _GEN_8275;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_30 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_30 <= _GEN_2592;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_30 <= _GEN_8276;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_31 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_31 <= _GEN_2593;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_31 <= _GEN_8277;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_32 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_32 <= _GEN_2594;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_32 <= _GEN_8278;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_33 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_33 <= _GEN_2595;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_33 <= _GEN_8279;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_34 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_34 <= _GEN_2596;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_34 <= _GEN_8280;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_35 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_35 <= _GEN_2597;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_35 <= _GEN_8281;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_36 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_36 <= _GEN_2598;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_36 <= _GEN_8282;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_37 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_37 <= _GEN_2599;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_37 <= _GEN_8283;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_38 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_38 <= _GEN_2600;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_38 <= _GEN_8284;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_39 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_39 <= _GEN_2601;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_39 <= _GEN_8285;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_40 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_40 <= _GEN_2602;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_40 <= _GEN_8286;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_41 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_41 <= _GEN_2603;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_41 <= _GEN_8287;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_42 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_42 <= _GEN_2604;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_42 <= _GEN_8288;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_43 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_43 <= _GEN_2605;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_43 <= _GEN_8289;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_44 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_44 <= _GEN_2606;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_44 <= _GEN_8290;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_45 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_45 <= _GEN_2607;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_45 <= _GEN_8291;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_46 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_46 <= _GEN_2608;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_46 <= _GEN_8292;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_47 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_47 <= _GEN_2609;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_47 <= _GEN_8293;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_48 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_48 <= _GEN_2610;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_48 <= _GEN_8294;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_49 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_49 <= _GEN_2611;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_49 <= _GEN_8295;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_50 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_50 <= _GEN_2612;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_50 <= _GEN_8296;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_51 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_51 <= _GEN_2613;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_51 <= _GEN_8297;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_52 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_52 <= _GEN_2614;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_52 <= _GEN_8298;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_53 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_53 <= _GEN_2615;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_53 <= _GEN_8299;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_54 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_54 <= _GEN_2616;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_54 <= _GEN_8300;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_55 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_55 <= _GEN_2617;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_55 <= _GEN_8301;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_56 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_56 <= _GEN_2618;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_56 <= _GEN_8302;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_57 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_57 <= _GEN_2619;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_57 <= _GEN_8303;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_58 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_58 <= _GEN_2620;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_58 <= _GEN_8304;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_59 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_59 <= _GEN_2621;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_59 <= _GEN_8305;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_60 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_60 <= _GEN_2622;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_60 <= _GEN_8306;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_61 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_61 <= _GEN_2623;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_61 <= _GEN_8307;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_62 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_62 <= _GEN_2624;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_62 <= _GEN_8308;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_63 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_63 <= _GEN_2625;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_63 <= _GEN_8309;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_64 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_64 <= _GEN_2626;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_64 <= _GEN_8310;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_65 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_65 <= _GEN_2627;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_65 <= _GEN_8311;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_66 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_66 <= _GEN_2628;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_66 <= _GEN_8312;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_67 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_67 <= _GEN_2629;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_67 <= _GEN_8313;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_68 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_68 <= _GEN_2630;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_68 <= _GEN_8314;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_69 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_69 <= _GEN_2631;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_69 <= _GEN_8315;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_70 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_70 <= _GEN_2632;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_70 <= _GEN_8316;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_71 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_71 <= _GEN_2633;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_71 <= _GEN_8317;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_72 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_72 <= _GEN_2634;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_72 <= _GEN_8318;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_73 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_73 <= _GEN_2635;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_73 <= _GEN_8319;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_74 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_74 <= _GEN_2636;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_74 <= _GEN_8320;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_75 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_75 <= _GEN_2637;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_75 <= _GEN_8321;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_76 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_76 <= _GEN_2638;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_76 <= _GEN_8322;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_77 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_77 <= _GEN_2639;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_77 <= _GEN_8323;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_78 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_78 <= _GEN_2640;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_78 <= _GEN_8324;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_79 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_79 <= _GEN_2641;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_79 <= _GEN_8325;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_80 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_80 <= _GEN_2642;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_80 <= _GEN_8326;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_81 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_81 <= _GEN_2643;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_81 <= _GEN_8327;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_82 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_82 <= _GEN_2644;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_82 <= _GEN_8328;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_83 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_83 <= _GEN_2645;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_83 <= _GEN_8329;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_84 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_84 <= _GEN_2646;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_84 <= _GEN_8330;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_85 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_85 <= _GEN_2647;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_85 <= _GEN_8331;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_86 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_86 <= _GEN_2648;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_86 <= _GEN_8332;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_87 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_87 <= _GEN_2649;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_87 <= _GEN_8333;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_88 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_88 <= _GEN_2650;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_88 <= _GEN_8334;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_89 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_89 <= _GEN_2651;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_89 <= _GEN_8335;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_90 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_90 <= _GEN_2652;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_90 <= _GEN_8336;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_91 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_91 <= _GEN_2653;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_91 <= _GEN_8337;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_92 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_92 <= _GEN_2654;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_92 <= _GEN_8338;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_93 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_93 <= _GEN_2655;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_93 <= _GEN_8339;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_94 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_94 <= _GEN_2656;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_94 <= _GEN_8340;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_95 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_95 <= _GEN_2657;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_95 <= _GEN_8341;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_96 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_96 <= _GEN_2658;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_96 <= _GEN_8342;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_97 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_97 <= _GEN_2659;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_97 <= _GEN_8343;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_98 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_98 <= _GEN_2660;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_98 <= _GEN_8344;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_99 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_99 <= _GEN_2661;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_99 <= _GEN_8345;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_100 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_100 <= _GEN_2662;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_100 <= _GEN_8346;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_101 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_101 <= _GEN_2663;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_101 <= _GEN_8347;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_102 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_102 <= _GEN_2664;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_102 <= _GEN_8348;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_103 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_103 <= _GEN_2665;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_103 <= _GEN_8349;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_104 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_104 <= _GEN_2666;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_104 <= _GEN_8350;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_105 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_105 <= _GEN_2667;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_105 <= _GEN_8351;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_106 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_106 <= _GEN_2668;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_106 <= _GEN_8352;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_107 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_107 <= _GEN_2669;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_107 <= _GEN_8353;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_108 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_108 <= _GEN_2670;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_108 <= _GEN_8354;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_109 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_109 <= _GEN_2671;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_109 <= _GEN_8355;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_110 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_110 <= _GEN_2672;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_110 <= _GEN_8356;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_111 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_111 <= _GEN_2673;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_111 <= _GEN_8357;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_112 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_112 <= _GEN_2674;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_112 <= _GEN_8358;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_113 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_113 <= _GEN_2675;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_113 <= _GEN_8359;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_114 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_114 <= _GEN_2676;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_114 <= _GEN_8360;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_115 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_115 <= _GEN_2677;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_115 <= _GEN_8361;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_116 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_116 <= _GEN_2678;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_116 <= _GEN_8362;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_117 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_117 <= _GEN_2679;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_117 <= _GEN_8363;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_118 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_118 <= _GEN_2680;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_118 <= _GEN_8364;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_119 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_119 <= _GEN_2681;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_119 <= _GEN_8365;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_120 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_120 <= _GEN_2682;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_120 <= _GEN_8366;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_121 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_121 <= _GEN_2683;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_121 <= _GEN_8367;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_122 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_122 <= _GEN_2684;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_122 <= _GEN_8368;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_123 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_123 <= _GEN_2685;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_123 <= _GEN_8369;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_124 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_124 <= _GEN_2686;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_124 <= _GEN_8370;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_125 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_125 <= _GEN_2687;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_125 <= _GEN_8371;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_126 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_126 <= _GEN_2688;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_126 <= _GEN_8372;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_127 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_127 <= _GEN_2689;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_127 <= _GEN_8373;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_128 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_128 <= _GEN_2690;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_128 <= _GEN_8374;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_129 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_129 <= _GEN_2691;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_129 <= _GEN_8375;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_130 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_130 <= _GEN_2692;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_130 <= _GEN_8376;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_131 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_131 <= _GEN_2693;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_131 <= _GEN_8377;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_132 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_132 <= _GEN_2694;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_132 <= _GEN_8378;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_133 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_133 <= _GEN_2695;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_133 <= _GEN_8379;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_134 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_134 <= _GEN_2696;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_134 <= _GEN_8380;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_135 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_135 <= _GEN_2697;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_135 <= _GEN_8381;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_136 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_136 <= _GEN_2698;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_136 <= _GEN_8382;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_137 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_137 <= _GEN_2699;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_137 <= _GEN_8383;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_138 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_138 <= _GEN_2700;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_138 <= _GEN_8384;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_139 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_139 <= _GEN_2701;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_139 <= _GEN_8385;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_140 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_140 <= _GEN_2702;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_140 <= _GEN_8386;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_141 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_141 <= _GEN_2703;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_141 <= _GEN_8387;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_142 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_142 <= _GEN_2704;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_142 <= _GEN_8388;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_143 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_143 <= _GEN_2705;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_143 <= _GEN_8389;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_144 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_144 <= _GEN_2706;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_144 <= _GEN_8390;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_145 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_145 <= _GEN_2707;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_145 <= _GEN_8391;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_146 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_146 <= _GEN_2708;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_146 <= _GEN_8392;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_147 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_147 <= _GEN_2709;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_147 <= _GEN_8393;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_148 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_148 <= _GEN_2710;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_148 <= _GEN_8394;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_149 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_149 <= _GEN_2711;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_149 <= _GEN_8395;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_150 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_150 <= _GEN_2712;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_150 <= _GEN_8396;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_151 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_151 <= _GEN_2713;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_151 <= _GEN_8397;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_152 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_152 <= _GEN_2714;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_152 <= _GEN_8398;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_153 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_153 <= _GEN_2715;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_153 <= _GEN_8399;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_154 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_154 <= _GEN_2716;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_154 <= _GEN_8400;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_155 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_155 <= _GEN_2717;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_155 <= _GEN_8401;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_156 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_156 <= _GEN_2718;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_156 <= _GEN_8402;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_157 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_157 <= _GEN_2719;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_157 <= _GEN_8403;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_158 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_158 <= _GEN_2720;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_158 <= _GEN_8404;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_159 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_159 <= _GEN_2721;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_159 <= _GEN_8405;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_160 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_160 <= _GEN_2722;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_160 <= _GEN_8406;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_161 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_161 <= _GEN_2723;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_161 <= _GEN_8407;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_162 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_162 <= _GEN_2724;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_162 <= _GEN_8408;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_163 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_163 <= _GEN_2725;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_163 <= _GEN_8409;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_164 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_164 <= _GEN_2726;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_164 <= _GEN_8410;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_165 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_165 <= _GEN_2727;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_165 <= _GEN_8411;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_166 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_166 <= _GEN_2728;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_166 <= _GEN_8412;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_167 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_167 <= _GEN_2729;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_167 <= _GEN_8413;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_168 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_168 <= _GEN_2730;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_168 <= _GEN_8414;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_169 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_169 <= _GEN_2731;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_169 <= _GEN_8415;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_170 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_170 <= _GEN_2732;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_170 <= _GEN_8416;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_171 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_171 <= _GEN_2733;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_171 <= _GEN_8417;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_172 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_172 <= _GEN_2734;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_172 <= _GEN_8418;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_173 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_173 <= _GEN_2735;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_173 <= _GEN_8419;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_174 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_174 <= _GEN_2736;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_174 <= _GEN_8420;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_175 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_175 <= _GEN_2737;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_175 <= _GEN_8421;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_176 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_176 <= _GEN_2738;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_176 <= _GEN_8422;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_177 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_177 <= _GEN_2739;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_177 <= _GEN_8423;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_178 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_178 <= _GEN_2740;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_178 <= _GEN_8424;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_179 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_179 <= _GEN_2741;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_179 <= _GEN_8425;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_180 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_180 <= _GEN_2742;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_180 <= _GEN_8426;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_181 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_181 <= _GEN_2743;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_181 <= _GEN_8427;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_182 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_182 <= _GEN_2744;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_182 <= _GEN_8428;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_183 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_183 <= _GEN_2745;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_183 <= _GEN_8429;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_184 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_184 <= _GEN_2746;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_184 <= _GEN_8430;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_185 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_185 <= _GEN_2747;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_185 <= _GEN_8431;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_186 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_186 <= _GEN_2748;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_186 <= _GEN_8432;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_187 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_187 <= _GEN_2749;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_187 <= _GEN_8433;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_188 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_188 <= _GEN_2750;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_188 <= _GEN_8434;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_189 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_189 <= _GEN_2751;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_189 <= _GEN_8435;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_190 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_190 <= _GEN_2752;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_190 <= _GEN_8436;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_191 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_191 <= _GEN_2753;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_191 <= _GEN_8437;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_192 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_192 <= _GEN_2754;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_192 <= _GEN_8438;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_193 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_193 <= _GEN_2755;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_193 <= _GEN_8439;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_194 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_194 <= _GEN_2756;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_194 <= _GEN_8440;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_195 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_195 <= _GEN_2757;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_195 <= _GEN_8441;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_196 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_196 <= _GEN_2758;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_196 <= _GEN_8442;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_197 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_197 <= _GEN_2759;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_197 <= _GEN_8443;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_198 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_198 <= _GEN_2760;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_198 <= _GEN_8444;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_199 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_199 <= _GEN_2761;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_199 <= _GEN_8445;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_200 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_200 <= _GEN_2762;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_200 <= _GEN_8446;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_201 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_201 <= _GEN_2763;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_201 <= _GEN_8447;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_202 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_202 <= _GEN_2764;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_202 <= _GEN_8448;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_203 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_203 <= _GEN_2765;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_203 <= _GEN_8449;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_204 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_204 <= _GEN_2766;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_204 <= _GEN_8450;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_205 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_205 <= _GEN_2767;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_205 <= _GEN_8451;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_206 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_206 <= _GEN_2768;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_206 <= _GEN_8452;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_207 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_207 <= _GEN_2769;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_207 <= _GEN_8453;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_208 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_208 <= _GEN_2770;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_208 <= _GEN_8454;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_209 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_209 <= _GEN_2771;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_209 <= _GEN_8455;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_210 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_210 <= _GEN_2772;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_210 <= _GEN_8456;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_211 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_211 <= _GEN_2773;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_211 <= _GEN_8457;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_212 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_212 <= _GEN_2774;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_212 <= _GEN_8458;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_213 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_213 <= _GEN_2775;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_213 <= _GEN_8459;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_214 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_214 <= _GEN_2776;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_214 <= _GEN_8460;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_215 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_215 <= _GEN_2777;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_215 <= _GEN_8461;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_216 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_216 <= _GEN_2778;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_216 <= _GEN_8462;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_217 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_217 <= _GEN_2779;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_217 <= _GEN_8463;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_218 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_218 <= _GEN_2780;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_218 <= _GEN_8464;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_219 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_219 <= _GEN_2781;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_219 <= _GEN_8465;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_220 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_220 <= _GEN_2782;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_220 <= _GEN_8466;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_221 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_221 <= _GEN_2783;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_221 <= _GEN_8467;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_222 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_222 <= _GEN_2784;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_222 <= _GEN_8468;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_223 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_223 <= _GEN_2785;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_223 <= _GEN_8469;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_224 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_224 <= _GEN_2786;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_224 <= _GEN_8470;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_225 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_225 <= _GEN_2787;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_225 <= _GEN_8471;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_226 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_226 <= _GEN_2788;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_226 <= _GEN_8472;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_227 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_227 <= _GEN_2789;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_227 <= _GEN_8473;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_228 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_228 <= _GEN_2790;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_228 <= _GEN_8474;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_229 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_229 <= _GEN_2791;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_229 <= _GEN_8475;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_230 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_230 <= _GEN_2792;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_230 <= _GEN_8476;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_231 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_231 <= _GEN_2793;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_231 <= _GEN_8477;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_232 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_232 <= _GEN_2794;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_232 <= _GEN_8478;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_233 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_233 <= _GEN_2795;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_233 <= _GEN_8479;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_234 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_234 <= _GEN_2796;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_234 <= _GEN_8480;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_235 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_235 <= _GEN_2797;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_235 <= _GEN_8481;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_236 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_236 <= _GEN_2798;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_236 <= _GEN_8482;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_237 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_237 <= _GEN_2799;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_237 <= _GEN_8483;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_238 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_238 <= _GEN_2800;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_238 <= _GEN_8484;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_239 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_239 <= _GEN_2801;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_239 <= _GEN_8485;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_240 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_240 <= _GEN_2802;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_240 <= _GEN_8486;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_241 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_241 <= _GEN_2803;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_241 <= _GEN_8487;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_242 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_242 <= _GEN_2804;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_242 <= _GEN_8488;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_243 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_243 <= _GEN_2805;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_243 <= _GEN_8489;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_244 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_244 <= _GEN_2806;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_244 <= _GEN_8490;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_245 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_245 <= _GEN_2807;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_245 <= _GEN_8491;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_246 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_246 <= _GEN_2808;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_246 <= _GEN_8492;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_247 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_247 <= _GEN_2809;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_247 <= _GEN_8493;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_248 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_248 <= _GEN_2810;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_248 <= _GEN_8494;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_249 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_249 <= _GEN_2811;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_249 <= _GEN_8495;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_250 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_250 <= _GEN_2812;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_250 <= _GEN_8496;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_251 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_251 <= _GEN_2813;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_251 <= _GEN_8497;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_252 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_252 <= _GEN_2814;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_252 <= _GEN_8498;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_253 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_253 <= _GEN_2815;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_253 <= _GEN_8499;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_254 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_254 <= _GEN_2816;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_254 <= _GEN_8500;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_255 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          offset_255 <= _GEN_2817;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        offset_255 <= _GEN_8501;
      end
    end
    if (reset) begin // @[Dcache.scala 26:22]
      state <= 3'h0; // @[Dcache.scala 26:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_dmem_data_valid) begin // @[Dcache.scala 125:28]
        state <= 3'h1; // @[Dcache.scala 126:15]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (~io_dmem_data_valid) begin // @[Dcache.scala 131:29]
        state <= 3'h0; // @[Dcache.scala 132:15]
      end else begin
        state <= _GEN_3078;
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      state <= _GEN_4364;
    end else begin
      state <= _GEN_7466;
    end
    if (reset) begin // @[Dcache.scala 46:28]
      data_ready <= 1'h0; // @[Dcache.scala 46:28]
    end else if (_T) begin // @[Conditional.scala 40:58]
      data_ready <= 1'h0; // @[Dcache.scala 123:18]
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
        data_ready <= _GEN_2818;
      end
    end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
      data_ready <= _GEN_7477;
    end
    if (reset) begin // @[Dcache.scala 116:28]
      cache_fill <= 1'h0; // @[Dcache.scala 116:28]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_4)) begin // @[Conditional.scala 39:67]
          cache_fill <= _GEN_7473;
        end
      end
    end
    if (reset) begin // @[Dcache.scala 117:28]
      cache_wen <= 1'h0; // @[Dcache.scala 117:28]
    end else if (_T) begin // @[Conditional.scala 40:58]
      cache_wen <= 1'h0; // @[Dcache.scala 124:18]
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
        cache_wen <= _GEN_2819;
      end
    end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
      cache_wen <= _GEN_7474;
    end
    if (reset) begin // @[Dcache.scala 118:28]
      cache_wdata <= 128'h0; // @[Dcache.scala 118:28]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          cache_wdata <= _GEN_2820;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        cache_wdata <= _GEN_7475;
      end
    end
    if (reset) begin // @[Dcache.scala 119:28]
      cache_strb <= 128'h0; // @[Dcache.scala 119:28]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (!(~io_dmem_data_valid)) begin // @[Dcache.scala 131:29]
          cache_strb <= _GEN_2821;
        end
      end else if (!(_T_4)) begin // @[Conditional.scala 39:67]
        cache_strb <= _GEN_7476;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_0 = _RAND_0[19:0];
  _RAND_1 = {1{`RANDOM}};
  tag_1 = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  tag_2 = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  tag_3 = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  tag_4 = _RAND_4[19:0];
  _RAND_5 = {1{`RANDOM}};
  tag_5 = _RAND_5[19:0];
  _RAND_6 = {1{`RANDOM}};
  tag_6 = _RAND_6[19:0];
  _RAND_7 = {1{`RANDOM}};
  tag_7 = _RAND_7[19:0];
  _RAND_8 = {1{`RANDOM}};
  tag_8 = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  tag_9 = _RAND_9[19:0];
  _RAND_10 = {1{`RANDOM}};
  tag_10 = _RAND_10[19:0];
  _RAND_11 = {1{`RANDOM}};
  tag_11 = _RAND_11[19:0];
  _RAND_12 = {1{`RANDOM}};
  tag_12 = _RAND_12[19:0];
  _RAND_13 = {1{`RANDOM}};
  tag_13 = _RAND_13[19:0];
  _RAND_14 = {1{`RANDOM}};
  tag_14 = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  tag_15 = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  tag_16 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  tag_17 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  tag_18 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  tag_19 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  tag_20 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  tag_21 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  tag_22 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  tag_23 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  tag_24 = _RAND_24[19:0];
  _RAND_25 = {1{`RANDOM}};
  tag_25 = _RAND_25[19:0];
  _RAND_26 = {1{`RANDOM}};
  tag_26 = _RAND_26[19:0];
  _RAND_27 = {1{`RANDOM}};
  tag_27 = _RAND_27[19:0];
  _RAND_28 = {1{`RANDOM}};
  tag_28 = _RAND_28[19:0];
  _RAND_29 = {1{`RANDOM}};
  tag_29 = _RAND_29[19:0];
  _RAND_30 = {1{`RANDOM}};
  tag_30 = _RAND_30[19:0];
  _RAND_31 = {1{`RANDOM}};
  tag_31 = _RAND_31[19:0];
  _RAND_32 = {1{`RANDOM}};
  tag_32 = _RAND_32[19:0];
  _RAND_33 = {1{`RANDOM}};
  tag_33 = _RAND_33[19:0];
  _RAND_34 = {1{`RANDOM}};
  tag_34 = _RAND_34[19:0];
  _RAND_35 = {1{`RANDOM}};
  tag_35 = _RAND_35[19:0];
  _RAND_36 = {1{`RANDOM}};
  tag_36 = _RAND_36[19:0];
  _RAND_37 = {1{`RANDOM}};
  tag_37 = _RAND_37[19:0];
  _RAND_38 = {1{`RANDOM}};
  tag_38 = _RAND_38[19:0];
  _RAND_39 = {1{`RANDOM}};
  tag_39 = _RAND_39[19:0];
  _RAND_40 = {1{`RANDOM}};
  tag_40 = _RAND_40[19:0];
  _RAND_41 = {1{`RANDOM}};
  tag_41 = _RAND_41[19:0];
  _RAND_42 = {1{`RANDOM}};
  tag_42 = _RAND_42[19:0];
  _RAND_43 = {1{`RANDOM}};
  tag_43 = _RAND_43[19:0];
  _RAND_44 = {1{`RANDOM}};
  tag_44 = _RAND_44[19:0];
  _RAND_45 = {1{`RANDOM}};
  tag_45 = _RAND_45[19:0];
  _RAND_46 = {1{`RANDOM}};
  tag_46 = _RAND_46[19:0];
  _RAND_47 = {1{`RANDOM}};
  tag_47 = _RAND_47[19:0];
  _RAND_48 = {1{`RANDOM}};
  tag_48 = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  tag_49 = _RAND_49[19:0];
  _RAND_50 = {1{`RANDOM}};
  tag_50 = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  tag_51 = _RAND_51[19:0];
  _RAND_52 = {1{`RANDOM}};
  tag_52 = _RAND_52[19:0];
  _RAND_53 = {1{`RANDOM}};
  tag_53 = _RAND_53[19:0];
  _RAND_54 = {1{`RANDOM}};
  tag_54 = _RAND_54[19:0];
  _RAND_55 = {1{`RANDOM}};
  tag_55 = _RAND_55[19:0];
  _RAND_56 = {1{`RANDOM}};
  tag_56 = _RAND_56[19:0];
  _RAND_57 = {1{`RANDOM}};
  tag_57 = _RAND_57[19:0];
  _RAND_58 = {1{`RANDOM}};
  tag_58 = _RAND_58[19:0];
  _RAND_59 = {1{`RANDOM}};
  tag_59 = _RAND_59[19:0];
  _RAND_60 = {1{`RANDOM}};
  tag_60 = _RAND_60[19:0];
  _RAND_61 = {1{`RANDOM}};
  tag_61 = _RAND_61[19:0];
  _RAND_62 = {1{`RANDOM}};
  tag_62 = _RAND_62[19:0];
  _RAND_63 = {1{`RANDOM}};
  tag_63 = _RAND_63[19:0];
  _RAND_64 = {1{`RANDOM}};
  tag_64 = _RAND_64[19:0];
  _RAND_65 = {1{`RANDOM}};
  tag_65 = _RAND_65[19:0];
  _RAND_66 = {1{`RANDOM}};
  tag_66 = _RAND_66[19:0];
  _RAND_67 = {1{`RANDOM}};
  tag_67 = _RAND_67[19:0];
  _RAND_68 = {1{`RANDOM}};
  tag_68 = _RAND_68[19:0];
  _RAND_69 = {1{`RANDOM}};
  tag_69 = _RAND_69[19:0];
  _RAND_70 = {1{`RANDOM}};
  tag_70 = _RAND_70[19:0];
  _RAND_71 = {1{`RANDOM}};
  tag_71 = _RAND_71[19:0];
  _RAND_72 = {1{`RANDOM}};
  tag_72 = _RAND_72[19:0];
  _RAND_73 = {1{`RANDOM}};
  tag_73 = _RAND_73[19:0];
  _RAND_74 = {1{`RANDOM}};
  tag_74 = _RAND_74[19:0];
  _RAND_75 = {1{`RANDOM}};
  tag_75 = _RAND_75[19:0];
  _RAND_76 = {1{`RANDOM}};
  tag_76 = _RAND_76[19:0];
  _RAND_77 = {1{`RANDOM}};
  tag_77 = _RAND_77[19:0];
  _RAND_78 = {1{`RANDOM}};
  tag_78 = _RAND_78[19:0];
  _RAND_79 = {1{`RANDOM}};
  tag_79 = _RAND_79[19:0];
  _RAND_80 = {1{`RANDOM}};
  tag_80 = _RAND_80[19:0];
  _RAND_81 = {1{`RANDOM}};
  tag_81 = _RAND_81[19:0];
  _RAND_82 = {1{`RANDOM}};
  tag_82 = _RAND_82[19:0];
  _RAND_83 = {1{`RANDOM}};
  tag_83 = _RAND_83[19:0];
  _RAND_84 = {1{`RANDOM}};
  tag_84 = _RAND_84[19:0];
  _RAND_85 = {1{`RANDOM}};
  tag_85 = _RAND_85[19:0];
  _RAND_86 = {1{`RANDOM}};
  tag_86 = _RAND_86[19:0];
  _RAND_87 = {1{`RANDOM}};
  tag_87 = _RAND_87[19:0];
  _RAND_88 = {1{`RANDOM}};
  tag_88 = _RAND_88[19:0];
  _RAND_89 = {1{`RANDOM}};
  tag_89 = _RAND_89[19:0];
  _RAND_90 = {1{`RANDOM}};
  tag_90 = _RAND_90[19:0];
  _RAND_91 = {1{`RANDOM}};
  tag_91 = _RAND_91[19:0];
  _RAND_92 = {1{`RANDOM}};
  tag_92 = _RAND_92[19:0];
  _RAND_93 = {1{`RANDOM}};
  tag_93 = _RAND_93[19:0];
  _RAND_94 = {1{`RANDOM}};
  tag_94 = _RAND_94[19:0];
  _RAND_95 = {1{`RANDOM}};
  tag_95 = _RAND_95[19:0];
  _RAND_96 = {1{`RANDOM}};
  tag_96 = _RAND_96[19:0];
  _RAND_97 = {1{`RANDOM}};
  tag_97 = _RAND_97[19:0];
  _RAND_98 = {1{`RANDOM}};
  tag_98 = _RAND_98[19:0];
  _RAND_99 = {1{`RANDOM}};
  tag_99 = _RAND_99[19:0];
  _RAND_100 = {1{`RANDOM}};
  tag_100 = _RAND_100[19:0];
  _RAND_101 = {1{`RANDOM}};
  tag_101 = _RAND_101[19:0];
  _RAND_102 = {1{`RANDOM}};
  tag_102 = _RAND_102[19:0];
  _RAND_103 = {1{`RANDOM}};
  tag_103 = _RAND_103[19:0];
  _RAND_104 = {1{`RANDOM}};
  tag_104 = _RAND_104[19:0];
  _RAND_105 = {1{`RANDOM}};
  tag_105 = _RAND_105[19:0];
  _RAND_106 = {1{`RANDOM}};
  tag_106 = _RAND_106[19:0];
  _RAND_107 = {1{`RANDOM}};
  tag_107 = _RAND_107[19:0];
  _RAND_108 = {1{`RANDOM}};
  tag_108 = _RAND_108[19:0];
  _RAND_109 = {1{`RANDOM}};
  tag_109 = _RAND_109[19:0];
  _RAND_110 = {1{`RANDOM}};
  tag_110 = _RAND_110[19:0];
  _RAND_111 = {1{`RANDOM}};
  tag_111 = _RAND_111[19:0];
  _RAND_112 = {1{`RANDOM}};
  tag_112 = _RAND_112[19:0];
  _RAND_113 = {1{`RANDOM}};
  tag_113 = _RAND_113[19:0];
  _RAND_114 = {1{`RANDOM}};
  tag_114 = _RAND_114[19:0];
  _RAND_115 = {1{`RANDOM}};
  tag_115 = _RAND_115[19:0];
  _RAND_116 = {1{`RANDOM}};
  tag_116 = _RAND_116[19:0];
  _RAND_117 = {1{`RANDOM}};
  tag_117 = _RAND_117[19:0];
  _RAND_118 = {1{`RANDOM}};
  tag_118 = _RAND_118[19:0];
  _RAND_119 = {1{`RANDOM}};
  tag_119 = _RAND_119[19:0];
  _RAND_120 = {1{`RANDOM}};
  tag_120 = _RAND_120[19:0];
  _RAND_121 = {1{`RANDOM}};
  tag_121 = _RAND_121[19:0];
  _RAND_122 = {1{`RANDOM}};
  tag_122 = _RAND_122[19:0];
  _RAND_123 = {1{`RANDOM}};
  tag_123 = _RAND_123[19:0];
  _RAND_124 = {1{`RANDOM}};
  tag_124 = _RAND_124[19:0];
  _RAND_125 = {1{`RANDOM}};
  tag_125 = _RAND_125[19:0];
  _RAND_126 = {1{`RANDOM}};
  tag_126 = _RAND_126[19:0];
  _RAND_127 = {1{`RANDOM}};
  tag_127 = _RAND_127[19:0];
  _RAND_128 = {1{`RANDOM}};
  tag_128 = _RAND_128[19:0];
  _RAND_129 = {1{`RANDOM}};
  tag_129 = _RAND_129[19:0];
  _RAND_130 = {1{`RANDOM}};
  tag_130 = _RAND_130[19:0];
  _RAND_131 = {1{`RANDOM}};
  tag_131 = _RAND_131[19:0];
  _RAND_132 = {1{`RANDOM}};
  tag_132 = _RAND_132[19:0];
  _RAND_133 = {1{`RANDOM}};
  tag_133 = _RAND_133[19:0];
  _RAND_134 = {1{`RANDOM}};
  tag_134 = _RAND_134[19:0];
  _RAND_135 = {1{`RANDOM}};
  tag_135 = _RAND_135[19:0];
  _RAND_136 = {1{`RANDOM}};
  tag_136 = _RAND_136[19:0];
  _RAND_137 = {1{`RANDOM}};
  tag_137 = _RAND_137[19:0];
  _RAND_138 = {1{`RANDOM}};
  tag_138 = _RAND_138[19:0];
  _RAND_139 = {1{`RANDOM}};
  tag_139 = _RAND_139[19:0];
  _RAND_140 = {1{`RANDOM}};
  tag_140 = _RAND_140[19:0];
  _RAND_141 = {1{`RANDOM}};
  tag_141 = _RAND_141[19:0];
  _RAND_142 = {1{`RANDOM}};
  tag_142 = _RAND_142[19:0];
  _RAND_143 = {1{`RANDOM}};
  tag_143 = _RAND_143[19:0];
  _RAND_144 = {1{`RANDOM}};
  tag_144 = _RAND_144[19:0];
  _RAND_145 = {1{`RANDOM}};
  tag_145 = _RAND_145[19:0];
  _RAND_146 = {1{`RANDOM}};
  tag_146 = _RAND_146[19:0];
  _RAND_147 = {1{`RANDOM}};
  tag_147 = _RAND_147[19:0];
  _RAND_148 = {1{`RANDOM}};
  tag_148 = _RAND_148[19:0];
  _RAND_149 = {1{`RANDOM}};
  tag_149 = _RAND_149[19:0];
  _RAND_150 = {1{`RANDOM}};
  tag_150 = _RAND_150[19:0];
  _RAND_151 = {1{`RANDOM}};
  tag_151 = _RAND_151[19:0];
  _RAND_152 = {1{`RANDOM}};
  tag_152 = _RAND_152[19:0];
  _RAND_153 = {1{`RANDOM}};
  tag_153 = _RAND_153[19:0];
  _RAND_154 = {1{`RANDOM}};
  tag_154 = _RAND_154[19:0];
  _RAND_155 = {1{`RANDOM}};
  tag_155 = _RAND_155[19:0];
  _RAND_156 = {1{`RANDOM}};
  tag_156 = _RAND_156[19:0];
  _RAND_157 = {1{`RANDOM}};
  tag_157 = _RAND_157[19:0];
  _RAND_158 = {1{`RANDOM}};
  tag_158 = _RAND_158[19:0];
  _RAND_159 = {1{`RANDOM}};
  tag_159 = _RAND_159[19:0];
  _RAND_160 = {1{`RANDOM}};
  tag_160 = _RAND_160[19:0];
  _RAND_161 = {1{`RANDOM}};
  tag_161 = _RAND_161[19:0];
  _RAND_162 = {1{`RANDOM}};
  tag_162 = _RAND_162[19:0];
  _RAND_163 = {1{`RANDOM}};
  tag_163 = _RAND_163[19:0];
  _RAND_164 = {1{`RANDOM}};
  tag_164 = _RAND_164[19:0];
  _RAND_165 = {1{`RANDOM}};
  tag_165 = _RAND_165[19:0];
  _RAND_166 = {1{`RANDOM}};
  tag_166 = _RAND_166[19:0];
  _RAND_167 = {1{`RANDOM}};
  tag_167 = _RAND_167[19:0];
  _RAND_168 = {1{`RANDOM}};
  tag_168 = _RAND_168[19:0];
  _RAND_169 = {1{`RANDOM}};
  tag_169 = _RAND_169[19:0];
  _RAND_170 = {1{`RANDOM}};
  tag_170 = _RAND_170[19:0];
  _RAND_171 = {1{`RANDOM}};
  tag_171 = _RAND_171[19:0];
  _RAND_172 = {1{`RANDOM}};
  tag_172 = _RAND_172[19:0];
  _RAND_173 = {1{`RANDOM}};
  tag_173 = _RAND_173[19:0];
  _RAND_174 = {1{`RANDOM}};
  tag_174 = _RAND_174[19:0];
  _RAND_175 = {1{`RANDOM}};
  tag_175 = _RAND_175[19:0];
  _RAND_176 = {1{`RANDOM}};
  tag_176 = _RAND_176[19:0];
  _RAND_177 = {1{`RANDOM}};
  tag_177 = _RAND_177[19:0];
  _RAND_178 = {1{`RANDOM}};
  tag_178 = _RAND_178[19:0];
  _RAND_179 = {1{`RANDOM}};
  tag_179 = _RAND_179[19:0];
  _RAND_180 = {1{`RANDOM}};
  tag_180 = _RAND_180[19:0];
  _RAND_181 = {1{`RANDOM}};
  tag_181 = _RAND_181[19:0];
  _RAND_182 = {1{`RANDOM}};
  tag_182 = _RAND_182[19:0];
  _RAND_183 = {1{`RANDOM}};
  tag_183 = _RAND_183[19:0];
  _RAND_184 = {1{`RANDOM}};
  tag_184 = _RAND_184[19:0];
  _RAND_185 = {1{`RANDOM}};
  tag_185 = _RAND_185[19:0];
  _RAND_186 = {1{`RANDOM}};
  tag_186 = _RAND_186[19:0];
  _RAND_187 = {1{`RANDOM}};
  tag_187 = _RAND_187[19:0];
  _RAND_188 = {1{`RANDOM}};
  tag_188 = _RAND_188[19:0];
  _RAND_189 = {1{`RANDOM}};
  tag_189 = _RAND_189[19:0];
  _RAND_190 = {1{`RANDOM}};
  tag_190 = _RAND_190[19:0];
  _RAND_191 = {1{`RANDOM}};
  tag_191 = _RAND_191[19:0];
  _RAND_192 = {1{`RANDOM}};
  tag_192 = _RAND_192[19:0];
  _RAND_193 = {1{`RANDOM}};
  tag_193 = _RAND_193[19:0];
  _RAND_194 = {1{`RANDOM}};
  tag_194 = _RAND_194[19:0];
  _RAND_195 = {1{`RANDOM}};
  tag_195 = _RAND_195[19:0];
  _RAND_196 = {1{`RANDOM}};
  tag_196 = _RAND_196[19:0];
  _RAND_197 = {1{`RANDOM}};
  tag_197 = _RAND_197[19:0];
  _RAND_198 = {1{`RANDOM}};
  tag_198 = _RAND_198[19:0];
  _RAND_199 = {1{`RANDOM}};
  tag_199 = _RAND_199[19:0];
  _RAND_200 = {1{`RANDOM}};
  tag_200 = _RAND_200[19:0];
  _RAND_201 = {1{`RANDOM}};
  tag_201 = _RAND_201[19:0];
  _RAND_202 = {1{`RANDOM}};
  tag_202 = _RAND_202[19:0];
  _RAND_203 = {1{`RANDOM}};
  tag_203 = _RAND_203[19:0];
  _RAND_204 = {1{`RANDOM}};
  tag_204 = _RAND_204[19:0];
  _RAND_205 = {1{`RANDOM}};
  tag_205 = _RAND_205[19:0];
  _RAND_206 = {1{`RANDOM}};
  tag_206 = _RAND_206[19:0];
  _RAND_207 = {1{`RANDOM}};
  tag_207 = _RAND_207[19:0];
  _RAND_208 = {1{`RANDOM}};
  tag_208 = _RAND_208[19:0];
  _RAND_209 = {1{`RANDOM}};
  tag_209 = _RAND_209[19:0];
  _RAND_210 = {1{`RANDOM}};
  tag_210 = _RAND_210[19:0];
  _RAND_211 = {1{`RANDOM}};
  tag_211 = _RAND_211[19:0];
  _RAND_212 = {1{`RANDOM}};
  tag_212 = _RAND_212[19:0];
  _RAND_213 = {1{`RANDOM}};
  tag_213 = _RAND_213[19:0];
  _RAND_214 = {1{`RANDOM}};
  tag_214 = _RAND_214[19:0];
  _RAND_215 = {1{`RANDOM}};
  tag_215 = _RAND_215[19:0];
  _RAND_216 = {1{`RANDOM}};
  tag_216 = _RAND_216[19:0];
  _RAND_217 = {1{`RANDOM}};
  tag_217 = _RAND_217[19:0];
  _RAND_218 = {1{`RANDOM}};
  tag_218 = _RAND_218[19:0];
  _RAND_219 = {1{`RANDOM}};
  tag_219 = _RAND_219[19:0];
  _RAND_220 = {1{`RANDOM}};
  tag_220 = _RAND_220[19:0];
  _RAND_221 = {1{`RANDOM}};
  tag_221 = _RAND_221[19:0];
  _RAND_222 = {1{`RANDOM}};
  tag_222 = _RAND_222[19:0];
  _RAND_223 = {1{`RANDOM}};
  tag_223 = _RAND_223[19:0];
  _RAND_224 = {1{`RANDOM}};
  tag_224 = _RAND_224[19:0];
  _RAND_225 = {1{`RANDOM}};
  tag_225 = _RAND_225[19:0];
  _RAND_226 = {1{`RANDOM}};
  tag_226 = _RAND_226[19:0];
  _RAND_227 = {1{`RANDOM}};
  tag_227 = _RAND_227[19:0];
  _RAND_228 = {1{`RANDOM}};
  tag_228 = _RAND_228[19:0];
  _RAND_229 = {1{`RANDOM}};
  tag_229 = _RAND_229[19:0];
  _RAND_230 = {1{`RANDOM}};
  tag_230 = _RAND_230[19:0];
  _RAND_231 = {1{`RANDOM}};
  tag_231 = _RAND_231[19:0];
  _RAND_232 = {1{`RANDOM}};
  tag_232 = _RAND_232[19:0];
  _RAND_233 = {1{`RANDOM}};
  tag_233 = _RAND_233[19:0];
  _RAND_234 = {1{`RANDOM}};
  tag_234 = _RAND_234[19:0];
  _RAND_235 = {1{`RANDOM}};
  tag_235 = _RAND_235[19:0];
  _RAND_236 = {1{`RANDOM}};
  tag_236 = _RAND_236[19:0];
  _RAND_237 = {1{`RANDOM}};
  tag_237 = _RAND_237[19:0];
  _RAND_238 = {1{`RANDOM}};
  tag_238 = _RAND_238[19:0];
  _RAND_239 = {1{`RANDOM}};
  tag_239 = _RAND_239[19:0];
  _RAND_240 = {1{`RANDOM}};
  tag_240 = _RAND_240[19:0];
  _RAND_241 = {1{`RANDOM}};
  tag_241 = _RAND_241[19:0];
  _RAND_242 = {1{`RANDOM}};
  tag_242 = _RAND_242[19:0];
  _RAND_243 = {1{`RANDOM}};
  tag_243 = _RAND_243[19:0];
  _RAND_244 = {1{`RANDOM}};
  tag_244 = _RAND_244[19:0];
  _RAND_245 = {1{`RANDOM}};
  tag_245 = _RAND_245[19:0];
  _RAND_246 = {1{`RANDOM}};
  tag_246 = _RAND_246[19:0];
  _RAND_247 = {1{`RANDOM}};
  tag_247 = _RAND_247[19:0];
  _RAND_248 = {1{`RANDOM}};
  tag_248 = _RAND_248[19:0];
  _RAND_249 = {1{`RANDOM}};
  tag_249 = _RAND_249[19:0];
  _RAND_250 = {1{`RANDOM}};
  tag_250 = _RAND_250[19:0];
  _RAND_251 = {1{`RANDOM}};
  tag_251 = _RAND_251[19:0];
  _RAND_252 = {1{`RANDOM}};
  tag_252 = _RAND_252[19:0];
  _RAND_253 = {1{`RANDOM}};
  tag_253 = _RAND_253[19:0];
  _RAND_254 = {1{`RANDOM}};
  tag_254 = _RAND_254[19:0];
  _RAND_255 = {1{`RANDOM}};
  tag_255 = _RAND_255[19:0];
  _RAND_256 = {1{`RANDOM}};
  valid_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_3 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_4 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_5 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_6 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_7 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_8 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_9 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_10 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_11 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_12 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_13 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_14 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_15 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_16 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_17 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_18 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_19 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_20 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_21 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_22 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_23 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_24 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_25 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_26 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_27 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_28 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_29 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_30 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_31 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_32 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_33 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_34 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_35 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_36 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_37 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_38 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_39 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_40 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_41 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_42 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_43 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_44 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_45 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_46 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_47 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_48 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_49 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_50 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_51 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_52 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_53 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_54 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_55 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_56 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_57 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_58 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_59 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_60 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_61 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_62 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_63 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_64 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_65 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_66 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_67 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid_68 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid_69 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid_70 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid_71 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid_72 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid_73 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid_74 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid_75 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid_76 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid_77 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid_78 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid_79 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid_80 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid_81 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid_82 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid_83 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid_84 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid_85 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid_86 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid_87 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid_88 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid_89 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid_90 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid_91 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid_92 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid_93 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid_94 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid_95 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid_96 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid_97 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid_98 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid_99 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid_100 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid_101 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid_102 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid_103 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid_104 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid_105 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid_106 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid_107 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid_108 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid_109 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid_110 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid_111 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid_112 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid_113 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid_114 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid_115 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid_116 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid_117 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid_118 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid_119 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid_120 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid_121 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid_122 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid_123 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid_124 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid_125 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid_126 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid_127 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  valid_128 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  valid_129 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  valid_130 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  valid_131 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  valid_132 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  valid_133 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  valid_134 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  valid_135 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  valid_136 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  valid_137 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  valid_138 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  valid_139 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  valid_140 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  valid_141 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  valid_142 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  valid_143 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  valid_144 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  valid_145 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  valid_146 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  valid_147 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  valid_148 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  valid_149 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  valid_150 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  valid_151 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  valid_152 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  valid_153 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  valid_154 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  valid_155 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  valid_156 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  valid_157 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  valid_158 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  valid_159 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  valid_160 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  valid_161 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  valid_162 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  valid_163 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  valid_164 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  valid_165 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  valid_166 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  valid_167 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  valid_168 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  valid_169 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  valid_170 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  valid_171 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  valid_172 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  valid_173 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  valid_174 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  valid_175 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  valid_176 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  valid_177 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  valid_178 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  valid_179 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  valid_180 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  valid_181 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  valid_182 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  valid_183 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  valid_184 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  valid_185 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  valid_186 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  valid_187 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  valid_188 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  valid_189 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  valid_190 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  valid_191 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  valid_192 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  valid_193 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  valid_194 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  valid_195 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  valid_196 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  valid_197 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  valid_198 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  valid_199 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  valid_200 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  valid_201 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  valid_202 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  valid_203 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  valid_204 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  valid_205 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  valid_206 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  valid_207 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  valid_208 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  valid_209 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  valid_210 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  valid_211 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  valid_212 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  valid_213 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  valid_214 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  valid_215 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  valid_216 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  valid_217 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  valid_218 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  valid_219 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  valid_220 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  valid_221 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  valid_222 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  valid_223 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  valid_224 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  valid_225 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  valid_226 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  valid_227 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  valid_228 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  valid_229 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  valid_230 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  valid_231 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  valid_232 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  valid_233 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  valid_234 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  valid_235 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  valid_236 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  valid_237 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  valid_238 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  valid_239 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  valid_240 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  valid_241 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  valid_242 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  valid_243 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  valid_244 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  valid_245 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  valid_246 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  valid_247 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  valid_248 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  valid_249 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  valid_250 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  valid_251 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  valid_252 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  valid_253 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  valid_254 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  valid_255 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  dirty_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  dirty_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  dirty_2 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  dirty_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  dirty_4 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  dirty_5 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  dirty_6 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  dirty_7 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  dirty_8 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  dirty_9 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  dirty_10 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  dirty_11 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  dirty_12 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  dirty_13 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  dirty_14 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  dirty_15 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  dirty_16 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  dirty_17 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  dirty_18 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  dirty_19 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  dirty_20 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  dirty_21 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  dirty_22 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  dirty_23 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  dirty_24 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  dirty_25 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  dirty_26 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  dirty_27 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  dirty_28 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  dirty_29 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  dirty_30 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  dirty_31 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  dirty_32 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  dirty_33 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  dirty_34 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  dirty_35 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  dirty_36 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  dirty_37 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  dirty_38 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  dirty_39 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  dirty_40 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  dirty_41 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  dirty_42 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  dirty_43 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  dirty_44 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  dirty_45 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  dirty_46 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  dirty_47 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  dirty_48 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  dirty_49 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  dirty_50 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  dirty_51 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  dirty_52 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  dirty_53 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  dirty_54 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  dirty_55 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  dirty_56 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  dirty_57 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  dirty_58 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  dirty_59 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  dirty_60 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  dirty_61 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  dirty_62 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  dirty_63 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  dirty_64 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  dirty_65 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  dirty_66 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  dirty_67 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  dirty_68 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  dirty_69 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  dirty_70 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  dirty_71 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  dirty_72 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  dirty_73 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  dirty_74 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  dirty_75 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  dirty_76 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  dirty_77 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  dirty_78 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  dirty_79 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  dirty_80 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  dirty_81 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  dirty_82 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  dirty_83 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  dirty_84 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  dirty_85 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  dirty_86 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  dirty_87 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  dirty_88 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  dirty_89 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  dirty_90 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  dirty_91 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  dirty_92 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  dirty_93 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  dirty_94 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  dirty_95 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  dirty_96 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  dirty_97 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  dirty_98 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  dirty_99 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  dirty_100 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  dirty_101 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  dirty_102 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  dirty_103 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  dirty_104 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  dirty_105 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  dirty_106 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  dirty_107 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  dirty_108 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  dirty_109 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  dirty_110 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  dirty_111 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  dirty_112 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  dirty_113 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  dirty_114 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  dirty_115 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  dirty_116 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  dirty_117 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  dirty_118 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  dirty_119 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  dirty_120 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  dirty_121 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  dirty_122 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  dirty_123 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  dirty_124 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  dirty_125 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  dirty_126 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  dirty_127 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  dirty_128 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  dirty_129 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  dirty_130 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  dirty_131 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  dirty_132 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  dirty_133 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  dirty_134 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  dirty_135 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  dirty_136 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  dirty_137 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  dirty_138 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  dirty_139 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  dirty_140 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  dirty_141 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  dirty_142 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  dirty_143 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  dirty_144 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  dirty_145 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  dirty_146 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  dirty_147 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  dirty_148 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  dirty_149 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  dirty_150 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  dirty_151 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  dirty_152 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  dirty_153 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  dirty_154 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  dirty_155 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  dirty_156 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  dirty_157 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  dirty_158 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  dirty_159 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  dirty_160 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  dirty_161 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  dirty_162 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  dirty_163 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  dirty_164 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  dirty_165 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  dirty_166 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  dirty_167 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  dirty_168 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  dirty_169 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  dirty_170 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  dirty_171 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  dirty_172 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  dirty_173 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  dirty_174 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  dirty_175 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  dirty_176 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  dirty_177 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  dirty_178 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  dirty_179 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  dirty_180 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  dirty_181 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  dirty_182 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  dirty_183 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  dirty_184 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  dirty_185 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  dirty_186 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  dirty_187 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  dirty_188 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  dirty_189 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  dirty_190 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  dirty_191 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  dirty_192 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  dirty_193 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  dirty_194 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  dirty_195 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  dirty_196 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  dirty_197 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  dirty_198 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  dirty_199 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  dirty_200 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  dirty_201 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  dirty_202 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  dirty_203 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  dirty_204 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  dirty_205 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  dirty_206 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  dirty_207 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  dirty_208 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  dirty_209 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  dirty_210 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  dirty_211 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  dirty_212 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  dirty_213 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  dirty_214 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  dirty_215 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  dirty_216 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  dirty_217 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  dirty_218 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  dirty_219 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  dirty_220 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  dirty_221 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  dirty_222 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  dirty_223 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  dirty_224 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  dirty_225 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  dirty_226 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  dirty_227 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  dirty_228 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  dirty_229 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  dirty_230 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  dirty_231 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  dirty_232 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  dirty_233 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  dirty_234 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  dirty_235 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  dirty_236 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  dirty_237 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  dirty_238 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  dirty_239 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  dirty_240 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  dirty_241 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  dirty_242 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  dirty_243 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  dirty_244 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  dirty_245 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  dirty_246 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  dirty_247 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  dirty_248 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  dirty_249 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  dirty_250 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  dirty_251 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  dirty_252 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  dirty_253 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  dirty_254 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  dirty_255 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  offset_0 = _RAND_768[3:0];
  _RAND_769 = {1{`RANDOM}};
  offset_1 = _RAND_769[3:0];
  _RAND_770 = {1{`RANDOM}};
  offset_2 = _RAND_770[3:0];
  _RAND_771 = {1{`RANDOM}};
  offset_3 = _RAND_771[3:0];
  _RAND_772 = {1{`RANDOM}};
  offset_4 = _RAND_772[3:0];
  _RAND_773 = {1{`RANDOM}};
  offset_5 = _RAND_773[3:0];
  _RAND_774 = {1{`RANDOM}};
  offset_6 = _RAND_774[3:0];
  _RAND_775 = {1{`RANDOM}};
  offset_7 = _RAND_775[3:0];
  _RAND_776 = {1{`RANDOM}};
  offset_8 = _RAND_776[3:0];
  _RAND_777 = {1{`RANDOM}};
  offset_9 = _RAND_777[3:0];
  _RAND_778 = {1{`RANDOM}};
  offset_10 = _RAND_778[3:0];
  _RAND_779 = {1{`RANDOM}};
  offset_11 = _RAND_779[3:0];
  _RAND_780 = {1{`RANDOM}};
  offset_12 = _RAND_780[3:0];
  _RAND_781 = {1{`RANDOM}};
  offset_13 = _RAND_781[3:0];
  _RAND_782 = {1{`RANDOM}};
  offset_14 = _RAND_782[3:0];
  _RAND_783 = {1{`RANDOM}};
  offset_15 = _RAND_783[3:0];
  _RAND_784 = {1{`RANDOM}};
  offset_16 = _RAND_784[3:0];
  _RAND_785 = {1{`RANDOM}};
  offset_17 = _RAND_785[3:0];
  _RAND_786 = {1{`RANDOM}};
  offset_18 = _RAND_786[3:0];
  _RAND_787 = {1{`RANDOM}};
  offset_19 = _RAND_787[3:0];
  _RAND_788 = {1{`RANDOM}};
  offset_20 = _RAND_788[3:0];
  _RAND_789 = {1{`RANDOM}};
  offset_21 = _RAND_789[3:0];
  _RAND_790 = {1{`RANDOM}};
  offset_22 = _RAND_790[3:0];
  _RAND_791 = {1{`RANDOM}};
  offset_23 = _RAND_791[3:0];
  _RAND_792 = {1{`RANDOM}};
  offset_24 = _RAND_792[3:0];
  _RAND_793 = {1{`RANDOM}};
  offset_25 = _RAND_793[3:0];
  _RAND_794 = {1{`RANDOM}};
  offset_26 = _RAND_794[3:0];
  _RAND_795 = {1{`RANDOM}};
  offset_27 = _RAND_795[3:0];
  _RAND_796 = {1{`RANDOM}};
  offset_28 = _RAND_796[3:0];
  _RAND_797 = {1{`RANDOM}};
  offset_29 = _RAND_797[3:0];
  _RAND_798 = {1{`RANDOM}};
  offset_30 = _RAND_798[3:0];
  _RAND_799 = {1{`RANDOM}};
  offset_31 = _RAND_799[3:0];
  _RAND_800 = {1{`RANDOM}};
  offset_32 = _RAND_800[3:0];
  _RAND_801 = {1{`RANDOM}};
  offset_33 = _RAND_801[3:0];
  _RAND_802 = {1{`RANDOM}};
  offset_34 = _RAND_802[3:0];
  _RAND_803 = {1{`RANDOM}};
  offset_35 = _RAND_803[3:0];
  _RAND_804 = {1{`RANDOM}};
  offset_36 = _RAND_804[3:0];
  _RAND_805 = {1{`RANDOM}};
  offset_37 = _RAND_805[3:0];
  _RAND_806 = {1{`RANDOM}};
  offset_38 = _RAND_806[3:0];
  _RAND_807 = {1{`RANDOM}};
  offset_39 = _RAND_807[3:0];
  _RAND_808 = {1{`RANDOM}};
  offset_40 = _RAND_808[3:0];
  _RAND_809 = {1{`RANDOM}};
  offset_41 = _RAND_809[3:0];
  _RAND_810 = {1{`RANDOM}};
  offset_42 = _RAND_810[3:0];
  _RAND_811 = {1{`RANDOM}};
  offset_43 = _RAND_811[3:0];
  _RAND_812 = {1{`RANDOM}};
  offset_44 = _RAND_812[3:0];
  _RAND_813 = {1{`RANDOM}};
  offset_45 = _RAND_813[3:0];
  _RAND_814 = {1{`RANDOM}};
  offset_46 = _RAND_814[3:0];
  _RAND_815 = {1{`RANDOM}};
  offset_47 = _RAND_815[3:0];
  _RAND_816 = {1{`RANDOM}};
  offset_48 = _RAND_816[3:0];
  _RAND_817 = {1{`RANDOM}};
  offset_49 = _RAND_817[3:0];
  _RAND_818 = {1{`RANDOM}};
  offset_50 = _RAND_818[3:0];
  _RAND_819 = {1{`RANDOM}};
  offset_51 = _RAND_819[3:0];
  _RAND_820 = {1{`RANDOM}};
  offset_52 = _RAND_820[3:0];
  _RAND_821 = {1{`RANDOM}};
  offset_53 = _RAND_821[3:0];
  _RAND_822 = {1{`RANDOM}};
  offset_54 = _RAND_822[3:0];
  _RAND_823 = {1{`RANDOM}};
  offset_55 = _RAND_823[3:0];
  _RAND_824 = {1{`RANDOM}};
  offset_56 = _RAND_824[3:0];
  _RAND_825 = {1{`RANDOM}};
  offset_57 = _RAND_825[3:0];
  _RAND_826 = {1{`RANDOM}};
  offset_58 = _RAND_826[3:0];
  _RAND_827 = {1{`RANDOM}};
  offset_59 = _RAND_827[3:0];
  _RAND_828 = {1{`RANDOM}};
  offset_60 = _RAND_828[3:0];
  _RAND_829 = {1{`RANDOM}};
  offset_61 = _RAND_829[3:0];
  _RAND_830 = {1{`RANDOM}};
  offset_62 = _RAND_830[3:0];
  _RAND_831 = {1{`RANDOM}};
  offset_63 = _RAND_831[3:0];
  _RAND_832 = {1{`RANDOM}};
  offset_64 = _RAND_832[3:0];
  _RAND_833 = {1{`RANDOM}};
  offset_65 = _RAND_833[3:0];
  _RAND_834 = {1{`RANDOM}};
  offset_66 = _RAND_834[3:0];
  _RAND_835 = {1{`RANDOM}};
  offset_67 = _RAND_835[3:0];
  _RAND_836 = {1{`RANDOM}};
  offset_68 = _RAND_836[3:0];
  _RAND_837 = {1{`RANDOM}};
  offset_69 = _RAND_837[3:0];
  _RAND_838 = {1{`RANDOM}};
  offset_70 = _RAND_838[3:0];
  _RAND_839 = {1{`RANDOM}};
  offset_71 = _RAND_839[3:0];
  _RAND_840 = {1{`RANDOM}};
  offset_72 = _RAND_840[3:0];
  _RAND_841 = {1{`RANDOM}};
  offset_73 = _RAND_841[3:0];
  _RAND_842 = {1{`RANDOM}};
  offset_74 = _RAND_842[3:0];
  _RAND_843 = {1{`RANDOM}};
  offset_75 = _RAND_843[3:0];
  _RAND_844 = {1{`RANDOM}};
  offset_76 = _RAND_844[3:0];
  _RAND_845 = {1{`RANDOM}};
  offset_77 = _RAND_845[3:0];
  _RAND_846 = {1{`RANDOM}};
  offset_78 = _RAND_846[3:0];
  _RAND_847 = {1{`RANDOM}};
  offset_79 = _RAND_847[3:0];
  _RAND_848 = {1{`RANDOM}};
  offset_80 = _RAND_848[3:0];
  _RAND_849 = {1{`RANDOM}};
  offset_81 = _RAND_849[3:0];
  _RAND_850 = {1{`RANDOM}};
  offset_82 = _RAND_850[3:0];
  _RAND_851 = {1{`RANDOM}};
  offset_83 = _RAND_851[3:0];
  _RAND_852 = {1{`RANDOM}};
  offset_84 = _RAND_852[3:0];
  _RAND_853 = {1{`RANDOM}};
  offset_85 = _RAND_853[3:0];
  _RAND_854 = {1{`RANDOM}};
  offset_86 = _RAND_854[3:0];
  _RAND_855 = {1{`RANDOM}};
  offset_87 = _RAND_855[3:0];
  _RAND_856 = {1{`RANDOM}};
  offset_88 = _RAND_856[3:0];
  _RAND_857 = {1{`RANDOM}};
  offset_89 = _RAND_857[3:0];
  _RAND_858 = {1{`RANDOM}};
  offset_90 = _RAND_858[3:0];
  _RAND_859 = {1{`RANDOM}};
  offset_91 = _RAND_859[3:0];
  _RAND_860 = {1{`RANDOM}};
  offset_92 = _RAND_860[3:0];
  _RAND_861 = {1{`RANDOM}};
  offset_93 = _RAND_861[3:0];
  _RAND_862 = {1{`RANDOM}};
  offset_94 = _RAND_862[3:0];
  _RAND_863 = {1{`RANDOM}};
  offset_95 = _RAND_863[3:0];
  _RAND_864 = {1{`RANDOM}};
  offset_96 = _RAND_864[3:0];
  _RAND_865 = {1{`RANDOM}};
  offset_97 = _RAND_865[3:0];
  _RAND_866 = {1{`RANDOM}};
  offset_98 = _RAND_866[3:0];
  _RAND_867 = {1{`RANDOM}};
  offset_99 = _RAND_867[3:0];
  _RAND_868 = {1{`RANDOM}};
  offset_100 = _RAND_868[3:0];
  _RAND_869 = {1{`RANDOM}};
  offset_101 = _RAND_869[3:0];
  _RAND_870 = {1{`RANDOM}};
  offset_102 = _RAND_870[3:0];
  _RAND_871 = {1{`RANDOM}};
  offset_103 = _RAND_871[3:0];
  _RAND_872 = {1{`RANDOM}};
  offset_104 = _RAND_872[3:0];
  _RAND_873 = {1{`RANDOM}};
  offset_105 = _RAND_873[3:0];
  _RAND_874 = {1{`RANDOM}};
  offset_106 = _RAND_874[3:0];
  _RAND_875 = {1{`RANDOM}};
  offset_107 = _RAND_875[3:0];
  _RAND_876 = {1{`RANDOM}};
  offset_108 = _RAND_876[3:0];
  _RAND_877 = {1{`RANDOM}};
  offset_109 = _RAND_877[3:0];
  _RAND_878 = {1{`RANDOM}};
  offset_110 = _RAND_878[3:0];
  _RAND_879 = {1{`RANDOM}};
  offset_111 = _RAND_879[3:0];
  _RAND_880 = {1{`RANDOM}};
  offset_112 = _RAND_880[3:0];
  _RAND_881 = {1{`RANDOM}};
  offset_113 = _RAND_881[3:0];
  _RAND_882 = {1{`RANDOM}};
  offset_114 = _RAND_882[3:0];
  _RAND_883 = {1{`RANDOM}};
  offset_115 = _RAND_883[3:0];
  _RAND_884 = {1{`RANDOM}};
  offset_116 = _RAND_884[3:0];
  _RAND_885 = {1{`RANDOM}};
  offset_117 = _RAND_885[3:0];
  _RAND_886 = {1{`RANDOM}};
  offset_118 = _RAND_886[3:0];
  _RAND_887 = {1{`RANDOM}};
  offset_119 = _RAND_887[3:0];
  _RAND_888 = {1{`RANDOM}};
  offset_120 = _RAND_888[3:0];
  _RAND_889 = {1{`RANDOM}};
  offset_121 = _RAND_889[3:0];
  _RAND_890 = {1{`RANDOM}};
  offset_122 = _RAND_890[3:0];
  _RAND_891 = {1{`RANDOM}};
  offset_123 = _RAND_891[3:0];
  _RAND_892 = {1{`RANDOM}};
  offset_124 = _RAND_892[3:0];
  _RAND_893 = {1{`RANDOM}};
  offset_125 = _RAND_893[3:0];
  _RAND_894 = {1{`RANDOM}};
  offset_126 = _RAND_894[3:0];
  _RAND_895 = {1{`RANDOM}};
  offset_127 = _RAND_895[3:0];
  _RAND_896 = {1{`RANDOM}};
  offset_128 = _RAND_896[3:0];
  _RAND_897 = {1{`RANDOM}};
  offset_129 = _RAND_897[3:0];
  _RAND_898 = {1{`RANDOM}};
  offset_130 = _RAND_898[3:0];
  _RAND_899 = {1{`RANDOM}};
  offset_131 = _RAND_899[3:0];
  _RAND_900 = {1{`RANDOM}};
  offset_132 = _RAND_900[3:0];
  _RAND_901 = {1{`RANDOM}};
  offset_133 = _RAND_901[3:0];
  _RAND_902 = {1{`RANDOM}};
  offset_134 = _RAND_902[3:0];
  _RAND_903 = {1{`RANDOM}};
  offset_135 = _RAND_903[3:0];
  _RAND_904 = {1{`RANDOM}};
  offset_136 = _RAND_904[3:0];
  _RAND_905 = {1{`RANDOM}};
  offset_137 = _RAND_905[3:0];
  _RAND_906 = {1{`RANDOM}};
  offset_138 = _RAND_906[3:0];
  _RAND_907 = {1{`RANDOM}};
  offset_139 = _RAND_907[3:0];
  _RAND_908 = {1{`RANDOM}};
  offset_140 = _RAND_908[3:0];
  _RAND_909 = {1{`RANDOM}};
  offset_141 = _RAND_909[3:0];
  _RAND_910 = {1{`RANDOM}};
  offset_142 = _RAND_910[3:0];
  _RAND_911 = {1{`RANDOM}};
  offset_143 = _RAND_911[3:0];
  _RAND_912 = {1{`RANDOM}};
  offset_144 = _RAND_912[3:0];
  _RAND_913 = {1{`RANDOM}};
  offset_145 = _RAND_913[3:0];
  _RAND_914 = {1{`RANDOM}};
  offset_146 = _RAND_914[3:0];
  _RAND_915 = {1{`RANDOM}};
  offset_147 = _RAND_915[3:0];
  _RAND_916 = {1{`RANDOM}};
  offset_148 = _RAND_916[3:0];
  _RAND_917 = {1{`RANDOM}};
  offset_149 = _RAND_917[3:0];
  _RAND_918 = {1{`RANDOM}};
  offset_150 = _RAND_918[3:0];
  _RAND_919 = {1{`RANDOM}};
  offset_151 = _RAND_919[3:0];
  _RAND_920 = {1{`RANDOM}};
  offset_152 = _RAND_920[3:0];
  _RAND_921 = {1{`RANDOM}};
  offset_153 = _RAND_921[3:0];
  _RAND_922 = {1{`RANDOM}};
  offset_154 = _RAND_922[3:0];
  _RAND_923 = {1{`RANDOM}};
  offset_155 = _RAND_923[3:0];
  _RAND_924 = {1{`RANDOM}};
  offset_156 = _RAND_924[3:0];
  _RAND_925 = {1{`RANDOM}};
  offset_157 = _RAND_925[3:0];
  _RAND_926 = {1{`RANDOM}};
  offset_158 = _RAND_926[3:0];
  _RAND_927 = {1{`RANDOM}};
  offset_159 = _RAND_927[3:0];
  _RAND_928 = {1{`RANDOM}};
  offset_160 = _RAND_928[3:0];
  _RAND_929 = {1{`RANDOM}};
  offset_161 = _RAND_929[3:0];
  _RAND_930 = {1{`RANDOM}};
  offset_162 = _RAND_930[3:0];
  _RAND_931 = {1{`RANDOM}};
  offset_163 = _RAND_931[3:0];
  _RAND_932 = {1{`RANDOM}};
  offset_164 = _RAND_932[3:0];
  _RAND_933 = {1{`RANDOM}};
  offset_165 = _RAND_933[3:0];
  _RAND_934 = {1{`RANDOM}};
  offset_166 = _RAND_934[3:0];
  _RAND_935 = {1{`RANDOM}};
  offset_167 = _RAND_935[3:0];
  _RAND_936 = {1{`RANDOM}};
  offset_168 = _RAND_936[3:0];
  _RAND_937 = {1{`RANDOM}};
  offset_169 = _RAND_937[3:0];
  _RAND_938 = {1{`RANDOM}};
  offset_170 = _RAND_938[3:0];
  _RAND_939 = {1{`RANDOM}};
  offset_171 = _RAND_939[3:0];
  _RAND_940 = {1{`RANDOM}};
  offset_172 = _RAND_940[3:0];
  _RAND_941 = {1{`RANDOM}};
  offset_173 = _RAND_941[3:0];
  _RAND_942 = {1{`RANDOM}};
  offset_174 = _RAND_942[3:0];
  _RAND_943 = {1{`RANDOM}};
  offset_175 = _RAND_943[3:0];
  _RAND_944 = {1{`RANDOM}};
  offset_176 = _RAND_944[3:0];
  _RAND_945 = {1{`RANDOM}};
  offset_177 = _RAND_945[3:0];
  _RAND_946 = {1{`RANDOM}};
  offset_178 = _RAND_946[3:0];
  _RAND_947 = {1{`RANDOM}};
  offset_179 = _RAND_947[3:0];
  _RAND_948 = {1{`RANDOM}};
  offset_180 = _RAND_948[3:0];
  _RAND_949 = {1{`RANDOM}};
  offset_181 = _RAND_949[3:0];
  _RAND_950 = {1{`RANDOM}};
  offset_182 = _RAND_950[3:0];
  _RAND_951 = {1{`RANDOM}};
  offset_183 = _RAND_951[3:0];
  _RAND_952 = {1{`RANDOM}};
  offset_184 = _RAND_952[3:0];
  _RAND_953 = {1{`RANDOM}};
  offset_185 = _RAND_953[3:0];
  _RAND_954 = {1{`RANDOM}};
  offset_186 = _RAND_954[3:0];
  _RAND_955 = {1{`RANDOM}};
  offset_187 = _RAND_955[3:0];
  _RAND_956 = {1{`RANDOM}};
  offset_188 = _RAND_956[3:0];
  _RAND_957 = {1{`RANDOM}};
  offset_189 = _RAND_957[3:0];
  _RAND_958 = {1{`RANDOM}};
  offset_190 = _RAND_958[3:0];
  _RAND_959 = {1{`RANDOM}};
  offset_191 = _RAND_959[3:0];
  _RAND_960 = {1{`RANDOM}};
  offset_192 = _RAND_960[3:0];
  _RAND_961 = {1{`RANDOM}};
  offset_193 = _RAND_961[3:0];
  _RAND_962 = {1{`RANDOM}};
  offset_194 = _RAND_962[3:0];
  _RAND_963 = {1{`RANDOM}};
  offset_195 = _RAND_963[3:0];
  _RAND_964 = {1{`RANDOM}};
  offset_196 = _RAND_964[3:0];
  _RAND_965 = {1{`RANDOM}};
  offset_197 = _RAND_965[3:0];
  _RAND_966 = {1{`RANDOM}};
  offset_198 = _RAND_966[3:0];
  _RAND_967 = {1{`RANDOM}};
  offset_199 = _RAND_967[3:0];
  _RAND_968 = {1{`RANDOM}};
  offset_200 = _RAND_968[3:0];
  _RAND_969 = {1{`RANDOM}};
  offset_201 = _RAND_969[3:0];
  _RAND_970 = {1{`RANDOM}};
  offset_202 = _RAND_970[3:0];
  _RAND_971 = {1{`RANDOM}};
  offset_203 = _RAND_971[3:0];
  _RAND_972 = {1{`RANDOM}};
  offset_204 = _RAND_972[3:0];
  _RAND_973 = {1{`RANDOM}};
  offset_205 = _RAND_973[3:0];
  _RAND_974 = {1{`RANDOM}};
  offset_206 = _RAND_974[3:0];
  _RAND_975 = {1{`RANDOM}};
  offset_207 = _RAND_975[3:0];
  _RAND_976 = {1{`RANDOM}};
  offset_208 = _RAND_976[3:0];
  _RAND_977 = {1{`RANDOM}};
  offset_209 = _RAND_977[3:0];
  _RAND_978 = {1{`RANDOM}};
  offset_210 = _RAND_978[3:0];
  _RAND_979 = {1{`RANDOM}};
  offset_211 = _RAND_979[3:0];
  _RAND_980 = {1{`RANDOM}};
  offset_212 = _RAND_980[3:0];
  _RAND_981 = {1{`RANDOM}};
  offset_213 = _RAND_981[3:0];
  _RAND_982 = {1{`RANDOM}};
  offset_214 = _RAND_982[3:0];
  _RAND_983 = {1{`RANDOM}};
  offset_215 = _RAND_983[3:0];
  _RAND_984 = {1{`RANDOM}};
  offset_216 = _RAND_984[3:0];
  _RAND_985 = {1{`RANDOM}};
  offset_217 = _RAND_985[3:0];
  _RAND_986 = {1{`RANDOM}};
  offset_218 = _RAND_986[3:0];
  _RAND_987 = {1{`RANDOM}};
  offset_219 = _RAND_987[3:0];
  _RAND_988 = {1{`RANDOM}};
  offset_220 = _RAND_988[3:0];
  _RAND_989 = {1{`RANDOM}};
  offset_221 = _RAND_989[3:0];
  _RAND_990 = {1{`RANDOM}};
  offset_222 = _RAND_990[3:0];
  _RAND_991 = {1{`RANDOM}};
  offset_223 = _RAND_991[3:0];
  _RAND_992 = {1{`RANDOM}};
  offset_224 = _RAND_992[3:0];
  _RAND_993 = {1{`RANDOM}};
  offset_225 = _RAND_993[3:0];
  _RAND_994 = {1{`RANDOM}};
  offset_226 = _RAND_994[3:0];
  _RAND_995 = {1{`RANDOM}};
  offset_227 = _RAND_995[3:0];
  _RAND_996 = {1{`RANDOM}};
  offset_228 = _RAND_996[3:0];
  _RAND_997 = {1{`RANDOM}};
  offset_229 = _RAND_997[3:0];
  _RAND_998 = {1{`RANDOM}};
  offset_230 = _RAND_998[3:0];
  _RAND_999 = {1{`RANDOM}};
  offset_231 = _RAND_999[3:0];
  _RAND_1000 = {1{`RANDOM}};
  offset_232 = _RAND_1000[3:0];
  _RAND_1001 = {1{`RANDOM}};
  offset_233 = _RAND_1001[3:0];
  _RAND_1002 = {1{`RANDOM}};
  offset_234 = _RAND_1002[3:0];
  _RAND_1003 = {1{`RANDOM}};
  offset_235 = _RAND_1003[3:0];
  _RAND_1004 = {1{`RANDOM}};
  offset_236 = _RAND_1004[3:0];
  _RAND_1005 = {1{`RANDOM}};
  offset_237 = _RAND_1005[3:0];
  _RAND_1006 = {1{`RANDOM}};
  offset_238 = _RAND_1006[3:0];
  _RAND_1007 = {1{`RANDOM}};
  offset_239 = _RAND_1007[3:0];
  _RAND_1008 = {1{`RANDOM}};
  offset_240 = _RAND_1008[3:0];
  _RAND_1009 = {1{`RANDOM}};
  offset_241 = _RAND_1009[3:0];
  _RAND_1010 = {1{`RANDOM}};
  offset_242 = _RAND_1010[3:0];
  _RAND_1011 = {1{`RANDOM}};
  offset_243 = _RAND_1011[3:0];
  _RAND_1012 = {1{`RANDOM}};
  offset_244 = _RAND_1012[3:0];
  _RAND_1013 = {1{`RANDOM}};
  offset_245 = _RAND_1013[3:0];
  _RAND_1014 = {1{`RANDOM}};
  offset_246 = _RAND_1014[3:0];
  _RAND_1015 = {1{`RANDOM}};
  offset_247 = _RAND_1015[3:0];
  _RAND_1016 = {1{`RANDOM}};
  offset_248 = _RAND_1016[3:0];
  _RAND_1017 = {1{`RANDOM}};
  offset_249 = _RAND_1017[3:0];
  _RAND_1018 = {1{`RANDOM}};
  offset_250 = _RAND_1018[3:0];
  _RAND_1019 = {1{`RANDOM}};
  offset_251 = _RAND_1019[3:0];
  _RAND_1020 = {1{`RANDOM}};
  offset_252 = _RAND_1020[3:0];
  _RAND_1021 = {1{`RANDOM}};
  offset_253 = _RAND_1021[3:0];
  _RAND_1022 = {1{`RANDOM}};
  offset_254 = _RAND_1022[3:0];
  _RAND_1023 = {1{`RANDOM}};
  offset_255 = _RAND_1023[3:0];
  _RAND_1024 = {1{`RANDOM}};
  state = _RAND_1024[2:0];
  _RAND_1025 = {1{`RANDOM}};
  data_ready = _RAND_1025[0:0];
  _RAND_1026 = {1{`RANDOM}};
  cache_fill = _RAND_1026[0:0];
  _RAND_1027 = {1{`RANDOM}};
  cache_wen = _RAND_1027[0:0];
  _RAND_1028 = {4{`RANDOM}};
  cache_wdata = _RAND_1028[127:0];
  _RAND_1029 = {4{`RANDOM}};
  cache_strb = _RAND_1029[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AxiLite2Axi(
  input          clock,
  input          reset,
  input          io_out_aw_ready,
  output         io_out_aw_valid,
  output [31:0]  io_out_aw_bits_addr,
  input          io_out_w_ready,
  output         io_out_w_valid,
  output [63:0]  io_out_w_bits_data,
  output [7:0]   io_out_w_bits_strb,
  output         io_out_w_bits_last,
  output         io_out_b_ready,
  input          io_out_b_valid,
  input          io_out_ar_ready,
  output         io_out_ar_valid,
  output [31:0]  io_out_ar_bits_addr,
  output         io_out_r_ready,
  input          io_out_r_valid,
  input  [63:0]  io_out_r_bits_data,
  input          io_out_r_bits_last,
  input          io_imem_inst_valid,
  output         io_imem_inst_ready,
  input  [31:0]  io_imem_inst_addr,
  output [127:0] io_imem_inst_read,
  input          io_dmem_data_valid,
  output         io_dmem_data_ready,
  input          io_dmem_data_req,
  input  [31:0]  io_dmem_data_addr,
  input  [7:0]   io_dmem_data_strb,
  output [127:0] io_dmem_data_read,
  input  [127:0] io_dmem_data_write
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  data_ren = io_dmem_data_valid & ~io_dmem_data_req; // @[AXI.scala 123:30]
  wire  data_wen = io_dmem_data_valid & io_dmem_data_req; // @[AXI.scala 124:30]
  wire  aw_hs = io_out_aw_ready & io_out_aw_valid; // @[AXI.scala 126:33]
  wire  w_hs = io_out_w_ready & io_out_w_valid; // @[AXI.scala 127:33]
  wire  b_hs = io_out_b_ready & io_out_b_valid; // @[AXI.scala 128:33]
  wire  ar_hs = io_out_ar_ready & io_out_ar_valid; // @[AXI.scala 129:33]
  wire  r_hs = io_out_r_ready & io_out_r_valid; // @[AXI.scala 130:33]
  wire  w_done = w_hs & io_out_w_bits_last; // @[AXI.scala 132:25]
  wire  r_done = r_hs & io_out_r_bits_last; // @[AXI.scala 133:25]
  reg [2:0] r_state; // @[AXI.scala 136:24]
  reg [2:0] w_state; // @[AXI.scala 139:24]
  wire  _T = 3'h0 == r_state; // @[Conditional.scala 37:30]
  wire  _T_1 = 3'h1 == r_state; // @[Conditional.scala 37:30]
  wire  _T_2 = 3'h2 == r_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_3 = r_done ? 3'h3 : r_state; // @[AXI.scala 156:21 AXI.scala 157:17 AXI.scala 136:24]
  wire  _T_3 = 3'h3 == r_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_4 = data_ren ? 3'h4 : 3'h0; // @[AXI.scala 161:23 AXI.scala 162:17 AXI.scala 165:17]
  wire  _T_4 = 3'h4 == r_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_5 = ar_hs ? 3'h5 : r_state; // @[AXI.scala 169:20 AXI.scala 170:17 AXI.scala 136:24]
  wire  _T_5 = 3'h5 == r_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_6 = r_done ? 3'h6 : r_state; // @[AXI.scala 174:21 AXI.scala 175:17 AXI.scala 136:24]
  wire  _T_6 = 3'h6 == r_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_7 = _T_6 ? 3'h0 : r_state; // @[Conditional.scala 39:67 AXI.scala 179:15 AXI.scala 136:24]
  wire [2:0] _GEN_8 = _T_5 ? _GEN_6 : _GEN_7; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_9 = _T_4 ? _GEN_5 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_3 ? _GEN_4 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _T_7 = 3'h0 == w_state; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h1 == w_state; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h2 == w_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_16 = w_done ? 3'h3 : w_state; // @[AXI.scala 195:21 AXI.scala 196:17 AXI.scala 139:24]
  wire  _T_10 = 3'h3 == w_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_17 = b_hs ? 3'h4 : w_state; // @[AXI.scala 200:19 AXI.scala 201:17 AXI.scala 139:24]
  wire  _T_11 = 3'h4 == w_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_18 = _T_11 ? 3'h0 : w_state; // @[Conditional.scala 39:67 AXI.scala 205:15 AXI.scala 139:24]
  wire [2:0] _GEN_19 = _T_10 ? _GEN_17 : _GEN_18; // @[Conditional.scala 39:67]
  reg  data_ok; // @[AXI.scala 209:24]
  wire  _T_12 = w_state == 3'h4; // @[AXI.scala 210:29]
  wire  _GEN_23 = ~data_wen ? 1'h0 : data_ok; // @[AXI.scala 213:25 AXI.scala 214:13 AXI.scala 209:24]
  wire  _GEN_24 = data_wen & w_state == 3'h4 | _GEN_23; // @[AXI.scala 210:46 AXI.scala 211:13]
  wire  _axi_addr_T = r_state == 3'h1; // @[AXI.scala 217:31]
  wire [31:0] _axi_addr_T_1 = io_imem_inst_addr & 32'hfffffff0; // @[AXI.scala 217:62]
  wire  _axi_addr_T_2 = r_state == 3'h4; // @[AXI.scala 218:31]
  wire [31:0] _axi_addr_T_3 = io_dmem_data_addr & 32'hfffffff0; // @[AXI.scala 218:62]
  wire [31:0] _axi_addr_T_4 = r_state == 3'h4 ? _axi_addr_T_3 : 32'h0; // @[AXI.scala 218:22]
  wire [27:0] axi_waddr_hi = io_dmem_data_addr[31:4]; // @[AXI.scala 219:49]
  wire [31:0] _axi_waddr_T = {axi_waddr_hi,4'h8}; // @[Cat.scala 30:58]
  reg [63:0] inst_read_h; // @[AXI.scala 265:28]
  reg [63:0] inst_read_l; // @[AXI.scala 266:28]
  reg [63:0] data_read_h; // @[AXI.scala 267:28]
  reg [63:0] data_read_l; // @[AXI.scala 268:28]
  assign io_out_aw_valid = w_state == 3'h1; // @[AXI.scala 238:34]
  assign io_out_aw_bits_addr = data_ok ? _axi_waddr_T : _axi_addr_T_3; // @[AXI.scala 219:22]
  assign io_out_w_valid = w_state == 3'h2; // @[AXI.scala 251:34]
  assign io_out_w_bits_data = data_ok ? io_dmem_data_write[127:64] : io_dmem_data_write[63:0]; // @[AXI.scala 252:29]
  assign io_out_w_bits_strb = io_dmem_data_strb; // @[AXI.scala 253:23]
  assign io_out_w_bits_last = 1'h1; // @[AXI.scala 254:23]
  assign io_out_b_ready = 1'h1; // @[AXI.scala 256:23]
  assign io_out_ar_valid = _axi_addr_T | _axi_addr_T_2; // @[AXI.scala 222:50]
  assign io_out_ar_bits_addr = r_state == 3'h1 ? _axi_addr_T_1 : _axi_addr_T_4; // @[AXI.scala 217:22]
  assign io_out_r_ready = 1'h1; // @[AXI.scala 235:23]
  assign io_imem_inst_ready = r_state == 3'h3; // @[AXI.scala 262:29]
  assign io_imem_inst_read = {inst_read_h,inst_read_l}; // @[Cat.scala 30:58]
  assign io_dmem_data_ready = r_state == 3'h6 | _T_12 & data_ok; // @[AXI.scala 263:45]
  assign io_dmem_data_read = {data_read_h,data_read_l}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if (reset) begin // @[AXI.scala 136:24]
      r_state <= 3'h0; // @[AXI.scala 136:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_imem_inst_valid) begin // @[AXI.scala 143:23]
        r_state <= 3'h1; // @[AXI.scala 144:17]
      end else if (data_ren) begin // @[AXI.scala 146:28]
        r_state <= 3'h4; // @[AXI.scala 147:17]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (ar_hs) begin // @[AXI.scala 151:20]
        r_state <= 3'h2; // @[AXI.scala 152:17]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      r_state <= _GEN_3;
    end else begin
      r_state <= _GEN_10;
    end
    if (reset) begin // @[AXI.scala 139:24]
      w_state <= 3'h0; // @[AXI.scala 139:24]
    end else if (_T_7) begin // @[Conditional.scala 40:58]
      if (data_wen) begin // @[AXI.scala 185:23]
        w_state <= 3'h1; // @[AXI.scala 186:17]
      end
    end else if (_T_8) begin // @[Conditional.scala 39:67]
      if (aw_hs) begin // @[AXI.scala 190:20]
        w_state <= 3'h2; // @[AXI.scala 191:17]
      end
    end else if (_T_9) begin // @[Conditional.scala 39:67]
      w_state <= _GEN_16;
    end else begin
      w_state <= _GEN_19;
    end
    if (reset) begin // @[AXI.scala 209:24]
      data_ok <= 1'h0; // @[AXI.scala 209:24]
    end else begin
      data_ok <= _GEN_24;
    end
    if (reset) begin // @[AXI.scala 265:28]
      inst_read_h <= 64'h0; // @[AXI.scala 265:28]
    end else if (r_hs) begin // @[AXI.scala 270:15]
      if (io_out_r_bits_last) begin // @[AXI.scala 271:28]
        inst_read_h <= io_out_r_bits_data; // @[AXI.scala 272:19]
      end
    end
    if (reset) begin // @[AXI.scala 266:28]
      inst_read_l <= 64'h0; // @[AXI.scala 266:28]
    end else if (r_hs) begin // @[AXI.scala 270:15]
      if (!(io_out_r_bits_last)) begin // @[AXI.scala 271:28]
        inst_read_l <= io_out_r_bits_data; // @[AXI.scala 276:19]
      end
    end
    if (reset) begin // @[AXI.scala 267:28]
      data_read_h <= 64'h0; // @[AXI.scala 267:28]
    end else if (r_hs) begin // @[AXI.scala 270:15]
      if (io_out_r_bits_last) begin // @[AXI.scala 271:28]
        data_read_h <= io_out_r_bits_data; // @[AXI.scala 273:19]
      end
    end
    if (reset) begin // @[AXI.scala 268:28]
      data_read_l <= 64'h0; // @[AXI.scala 268:28]
    end else if (r_hs) begin // @[AXI.scala 270:15]
      if (!(io_out_r_bits_last)) begin // @[AXI.scala 271:28]
        data_read_l <= io_out_r_bits_data; // @[AXI.scala 277:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  w_state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  data_ok = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  inst_read_h = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  inst_read_l = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  data_read_h = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  data_read_l = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimTop(
  input         clock,
  input         reset,
  input  [63:0] io_logCtrl_log_begin,
  input  [63:0] io_logCtrl_log_end,
  input  [63:0] io_logCtrl_log_level,
  input         io_perfInfo_clean,
  input         io_perfInfo_dump,
  output        io_uart_out_valid,
  output [7:0]  io_uart_out_ch,
  output        io_uart_in_valid,
  input  [7:0]  io_uart_in_ch,
  input         io_memAXI_0_aw_ready,
  output        io_memAXI_0_aw_valid,
  output [31:0] io_memAXI_0_aw_bits_addr,
  output [2:0]  io_memAXI_0_aw_bits_prot,
  output [3:0]  io_memAXI_0_aw_bits_id,
  output        io_memAXI_0_aw_bits_user,
  output [7:0]  io_memAXI_0_aw_bits_len,
  output [2:0]  io_memAXI_0_aw_bits_size,
  output [1:0]  io_memAXI_0_aw_bits_burst,
  output        io_memAXI_0_aw_bits_lock,
  output [3:0]  io_memAXI_0_aw_bits_cache,
  output [3:0]  io_memAXI_0_aw_bits_qos,
  input         io_memAXI_0_w_ready,
  output        io_memAXI_0_w_valid,
  output [63:0] io_memAXI_0_w_bits_data,
  output [7:0]  io_memAXI_0_w_bits_strb,
  output        io_memAXI_0_w_bits_last,
  output        io_memAXI_0_b_ready,
  input         io_memAXI_0_b_valid,
  input  [1:0]  io_memAXI_0_b_bits_resp,
  input  [3:0]  io_memAXI_0_b_bits_id,
  input         io_memAXI_0_b_bits_user,
  input         io_memAXI_0_ar_ready,
  output        io_memAXI_0_ar_valid,
  output [31:0] io_memAXI_0_ar_bits_addr,
  output [2:0]  io_memAXI_0_ar_bits_prot,
  output [3:0]  io_memAXI_0_ar_bits_id,
  output        io_memAXI_0_ar_bits_user,
  output [7:0]  io_memAXI_0_ar_bits_len,
  output [2:0]  io_memAXI_0_ar_bits_size,
  output [1:0]  io_memAXI_0_ar_bits_burst,
  output        io_memAXI_0_ar_bits_lock,
  output [3:0]  io_memAXI_0_ar_bits_cache,
  output [3:0]  io_memAXI_0_ar_bits_qos,
  output        io_memAXI_0_r_ready,
  input         io_memAXI_0_r_valid,
  input  [1:0]  io_memAXI_0_r_bits_resp,
  input  [63:0] io_memAXI_0_r_bits_data,
  input  [3:0]  io_memAXI_0_r_bits_id,
  input         io_memAXI_0_r_bits_user,
  input         io_memAXI_0_r_bits_last
);
  wire  core_clock; // @[SimTop.scala 15:20]
  wire  core_reset; // @[SimTop.scala 15:20]
  wire  core_io_imem_inst_valid; // @[SimTop.scala 15:20]
  wire  core_io_imem_inst_ready; // @[SimTop.scala 15:20]
  wire [31:0] core_io_imem_inst_addr; // @[SimTop.scala 15:20]
  wire [31:0] core_io_imem_inst_read; // @[SimTop.scala 15:20]
  wire  core_io_dmem_data_valid; // @[SimTop.scala 15:20]
  wire  core_io_dmem_data_ready; // @[SimTop.scala 15:20]
  wire  core_io_dmem_data_req; // @[SimTop.scala 15:20]
  wire [31:0] core_io_dmem_data_addr; // @[SimTop.scala 15:20]
  wire [1:0] core_io_dmem_data_size; // @[SimTop.scala 15:20]
  wire [7:0] core_io_dmem_data_strb; // @[SimTop.scala 15:20]
  wire [63:0] core_io_dmem_data_read; // @[SimTop.scala 15:20]
  wire [63:0] core_io_dmem_data_write; // @[SimTop.scala 15:20]
  wire  core_io_br_stall; // @[SimTop.scala 15:20]
  wire  icache_clock; // @[SimTop.scala 16:22]
  wire  icache_reset; // @[SimTop.scala 16:22]
  wire  icache_io_imem_inst_valid; // @[SimTop.scala 16:22]
  wire  icache_io_imem_inst_ready; // @[SimTop.scala 16:22]
  wire [31:0] icache_io_imem_inst_addr; // @[SimTop.scala 16:22]
  wire [31:0] icache_io_imem_inst_read; // @[SimTop.scala 16:22]
  wire  icache_io_out_inst_valid; // @[SimTop.scala 16:22]
  wire  icache_io_out_inst_ready; // @[SimTop.scala 16:22]
  wire [31:0] icache_io_out_inst_addr; // @[SimTop.scala 16:22]
  wire [127:0] icache_io_out_inst_read; // @[SimTop.scala 16:22]
  wire  icache_io_br_stall; // @[SimTop.scala 16:22]
  wire  dcache_clock; // @[SimTop.scala 17:22]
  wire  dcache_reset; // @[SimTop.scala 17:22]
  wire  dcache_io_dmem_data_valid; // @[SimTop.scala 17:22]
  wire  dcache_io_dmem_data_ready; // @[SimTop.scala 17:22]
  wire  dcache_io_dmem_data_req; // @[SimTop.scala 17:22]
  wire [31:0] dcache_io_dmem_data_addr; // @[SimTop.scala 17:22]
  wire [1:0] dcache_io_dmem_data_size; // @[SimTop.scala 17:22]
  wire [7:0] dcache_io_dmem_data_strb; // @[SimTop.scala 17:22]
  wire [63:0] dcache_io_dmem_data_read; // @[SimTop.scala 17:22]
  wire [63:0] dcache_io_dmem_data_write; // @[SimTop.scala 17:22]
  wire  dcache_io_out_data_valid; // @[SimTop.scala 17:22]
  wire  dcache_io_out_data_ready; // @[SimTop.scala 17:22]
  wire  dcache_io_out_data_req; // @[SimTop.scala 17:22]
  wire [31:0] dcache_io_out_data_addr; // @[SimTop.scala 17:22]
  wire [7:0] dcache_io_out_data_strb; // @[SimTop.scala 17:22]
  wire [127:0] dcache_io_out_data_read; // @[SimTop.scala 17:22]
  wire [127:0] dcache_io_out_data_write; // @[SimTop.scala 17:22]
  wire  top_clock; // @[SimTop.scala 19:19]
  wire  top_reset; // @[SimTop.scala 19:19]
  wire  top_io_out_aw_ready; // @[SimTop.scala 19:19]
  wire  top_io_out_aw_valid; // @[SimTop.scala 19:19]
  wire [31:0] top_io_out_aw_bits_addr; // @[SimTop.scala 19:19]
  wire  top_io_out_w_ready; // @[SimTop.scala 19:19]
  wire  top_io_out_w_valid; // @[SimTop.scala 19:19]
  wire [63:0] top_io_out_w_bits_data; // @[SimTop.scala 19:19]
  wire [7:0] top_io_out_w_bits_strb; // @[SimTop.scala 19:19]
  wire  top_io_out_w_bits_last; // @[SimTop.scala 19:19]
  wire  top_io_out_b_ready; // @[SimTop.scala 19:19]
  wire  top_io_out_b_valid; // @[SimTop.scala 19:19]
  wire  top_io_out_ar_ready; // @[SimTop.scala 19:19]
  wire  top_io_out_ar_valid; // @[SimTop.scala 19:19]
  wire [31:0] top_io_out_ar_bits_addr; // @[SimTop.scala 19:19]
  wire  top_io_out_r_ready; // @[SimTop.scala 19:19]
  wire  top_io_out_r_valid; // @[SimTop.scala 19:19]
  wire [63:0] top_io_out_r_bits_data; // @[SimTop.scala 19:19]
  wire  top_io_out_r_bits_last; // @[SimTop.scala 19:19]
  wire  top_io_imem_inst_valid; // @[SimTop.scala 19:19]
  wire  top_io_imem_inst_ready; // @[SimTop.scala 19:19]
  wire [31:0] top_io_imem_inst_addr; // @[SimTop.scala 19:19]
  wire [127:0] top_io_imem_inst_read; // @[SimTop.scala 19:19]
  wire  top_io_dmem_data_valid; // @[SimTop.scala 19:19]
  wire  top_io_dmem_data_ready; // @[SimTop.scala 19:19]
  wire  top_io_dmem_data_req; // @[SimTop.scala 19:19]
  wire [31:0] top_io_dmem_data_addr; // @[SimTop.scala 19:19]
  wire [7:0] top_io_dmem_data_strb; // @[SimTop.scala 19:19]
  wire [127:0] top_io_dmem_data_read; // @[SimTop.scala 19:19]
  wire [127:0] top_io_dmem_data_write; // @[SimTop.scala 19:19]
  Core core ( // @[SimTop.scala 15:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_inst_valid(core_io_imem_inst_valid),
    .io_imem_inst_ready(core_io_imem_inst_ready),
    .io_imem_inst_addr(core_io_imem_inst_addr),
    .io_imem_inst_read(core_io_imem_inst_read),
    .io_dmem_data_valid(core_io_dmem_data_valid),
    .io_dmem_data_ready(core_io_dmem_data_ready),
    .io_dmem_data_req(core_io_dmem_data_req),
    .io_dmem_data_addr(core_io_dmem_data_addr),
    .io_dmem_data_size(core_io_dmem_data_size),
    .io_dmem_data_strb(core_io_dmem_data_strb),
    .io_dmem_data_read(core_io_dmem_data_read),
    .io_dmem_data_write(core_io_dmem_data_write),
    .io_br_stall(core_io_br_stall)
  );
  Icache icache ( // @[SimTop.scala 16:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_imem_inst_valid(icache_io_imem_inst_valid),
    .io_imem_inst_ready(icache_io_imem_inst_ready),
    .io_imem_inst_addr(icache_io_imem_inst_addr),
    .io_imem_inst_read(icache_io_imem_inst_read),
    .io_out_inst_valid(icache_io_out_inst_valid),
    .io_out_inst_ready(icache_io_out_inst_ready),
    .io_out_inst_addr(icache_io_out_inst_addr),
    .io_out_inst_read(icache_io_out_inst_read),
    .io_br_stall(icache_io_br_stall)
  );
  Dcache dcache ( // @[SimTop.scala 17:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_dmem_data_valid(dcache_io_dmem_data_valid),
    .io_dmem_data_ready(dcache_io_dmem_data_ready),
    .io_dmem_data_req(dcache_io_dmem_data_req),
    .io_dmem_data_addr(dcache_io_dmem_data_addr),
    .io_dmem_data_size(dcache_io_dmem_data_size),
    .io_dmem_data_strb(dcache_io_dmem_data_strb),
    .io_dmem_data_read(dcache_io_dmem_data_read),
    .io_dmem_data_write(dcache_io_dmem_data_write),
    .io_out_data_valid(dcache_io_out_data_valid),
    .io_out_data_ready(dcache_io_out_data_ready),
    .io_out_data_req(dcache_io_out_data_req),
    .io_out_data_addr(dcache_io_out_data_addr),
    .io_out_data_strb(dcache_io_out_data_strb),
    .io_out_data_read(dcache_io_out_data_read),
    .io_out_data_write(dcache_io_out_data_write)
  );
  AxiLite2Axi top ( // @[SimTop.scala 19:19]
    .clock(top_clock),
    .reset(top_reset),
    .io_out_aw_ready(top_io_out_aw_ready),
    .io_out_aw_valid(top_io_out_aw_valid),
    .io_out_aw_bits_addr(top_io_out_aw_bits_addr),
    .io_out_w_ready(top_io_out_w_ready),
    .io_out_w_valid(top_io_out_w_valid),
    .io_out_w_bits_data(top_io_out_w_bits_data),
    .io_out_w_bits_strb(top_io_out_w_bits_strb),
    .io_out_w_bits_last(top_io_out_w_bits_last),
    .io_out_b_ready(top_io_out_b_ready),
    .io_out_b_valid(top_io_out_b_valid),
    .io_out_ar_ready(top_io_out_ar_ready),
    .io_out_ar_valid(top_io_out_ar_valid),
    .io_out_ar_bits_addr(top_io_out_ar_bits_addr),
    .io_out_r_ready(top_io_out_r_ready),
    .io_out_r_valid(top_io_out_r_valid),
    .io_out_r_bits_data(top_io_out_r_bits_data),
    .io_out_r_bits_last(top_io_out_r_bits_last),
    .io_imem_inst_valid(top_io_imem_inst_valid),
    .io_imem_inst_ready(top_io_imem_inst_ready),
    .io_imem_inst_addr(top_io_imem_inst_addr),
    .io_imem_inst_read(top_io_imem_inst_read),
    .io_dmem_data_valid(top_io_dmem_data_valid),
    .io_dmem_data_ready(top_io_dmem_data_ready),
    .io_dmem_data_req(top_io_dmem_data_req),
    .io_dmem_data_addr(top_io_dmem_data_addr),
    .io_dmem_data_strb(top_io_dmem_data_strb),
    .io_dmem_data_read(top_io_dmem_data_read),
    .io_dmem_data_write(top_io_dmem_data_write)
  );
  assign io_uart_out_valid = 1'h0; // @[SimTop.scala 39:21]
  assign io_uart_out_ch = 8'h0; // @[SimTop.scala 40:18]
  assign io_uart_in_valid = 1'h0; // @[SimTop.scala 41:20]
  assign io_memAXI_0_aw_valid = top_io_out_aw_valid; // @[SimTop.scala 33:18]
  assign io_memAXI_0_aw_bits_addr = top_io_out_aw_bits_addr; // @[SimTop.scala 33:18]
  assign io_memAXI_0_aw_bits_prot = 3'h0; // @[SimTop.scala 33:18]
  assign io_memAXI_0_aw_bits_id = 4'h0; // @[SimTop.scala 33:18]
  assign io_memAXI_0_aw_bits_user = 1'h0; // @[SimTop.scala 33:18]
  assign io_memAXI_0_aw_bits_len = 8'h0; // @[SimTop.scala 33:18]
  assign io_memAXI_0_aw_bits_size = 3'h3; // @[SimTop.scala 33:18]
  assign io_memAXI_0_aw_bits_burst = 2'h1; // @[SimTop.scala 33:18]
  assign io_memAXI_0_aw_bits_lock = 1'h0; // @[SimTop.scala 33:18]
  assign io_memAXI_0_aw_bits_cache = 4'h2; // @[SimTop.scala 33:18]
  assign io_memAXI_0_aw_bits_qos = 4'h0; // @[SimTop.scala 33:18]
  assign io_memAXI_0_w_valid = top_io_out_w_valid; // @[SimTop.scala 34:18]
  assign io_memAXI_0_w_bits_data = top_io_out_w_bits_data; // @[SimTop.scala 34:18]
  assign io_memAXI_0_w_bits_strb = top_io_out_w_bits_strb; // @[SimTop.scala 34:18]
  assign io_memAXI_0_w_bits_last = 1'h1; // @[SimTop.scala 34:18]
  assign io_memAXI_0_b_ready = 1'h1; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_valid = top_io_out_ar_valid; // @[SimTop.scala 36:18]
  assign io_memAXI_0_ar_bits_addr = top_io_out_ar_bits_addr; // @[SimTop.scala 36:18]
  assign io_memAXI_0_ar_bits_prot = 3'h0; // @[SimTop.scala 36:18]
  assign io_memAXI_0_ar_bits_id = 4'h0; // @[SimTop.scala 36:18]
  assign io_memAXI_0_ar_bits_user = 1'h0; // @[SimTop.scala 36:18]
  assign io_memAXI_0_ar_bits_len = 8'h1; // @[SimTop.scala 36:18]
  assign io_memAXI_0_ar_bits_size = 3'h3; // @[SimTop.scala 36:18]
  assign io_memAXI_0_ar_bits_burst = 2'h1; // @[SimTop.scala 36:18]
  assign io_memAXI_0_ar_bits_lock = 1'h0; // @[SimTop.scala 36:18]
  assign io_memAXI_0_ar_bits_cache = 4'h2; // @[SimTop.scala 36:18]
  assign io_memAXI_0_ar_bits_qos = 4'h0; // @[SimTop.scala 36:18]
  assign io_memAXI_0_r_ready = 1'h1; // @[SimTop.scala 37:18]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_imem_inst_ready = icache_io_imem_inst_ready; // @[SimTop.scala 21:17]
  assign core_io_imem_inst_read = icache_io_imem_inst_read; // @[SimTop.scala 21:17]
  assign core_io_dmem_data_ready = dcache_io_dmem_data_ready; // @[SimTop.scala 23:17]
  assign core_io_dmem_data_read = dcache_io_dmem_data_read; // @[SimTop.scala 23:17]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_imem_inst_valid = core_io_imem_inst_valid; // @[SimTop.scala 21:17]
  assign icache_io_imem_inst_addr = core_io_imem_inst_addr; // @[SimTop.scala 21:17]
  assign icache_io_out_inst_ready = top_io_imem_inst_ready; // @[SimTop.scala 22:17]
  assign icache_io_out_inst_read = top_io_imem_inst_read; // @[SimTop.scala 22:17]
  assign icache_io_br_stall = core_io_br_stall; // @[SimTop.scala 26:25]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_dmem_data_valid = core_io_dmem_data_valid; // @[SimTop.scala 23:17]
  assign dcache_io_dmem_data_req = core_io_dmem_data_req; // @[SimTop.scala 23:17]
  assign dcache_io_dmem_data_addr = core_io_dmem_data_addr; // @[SimTop.scala 23:17]
  assign dcache_io_dmem_data_size = core_io_dmem_data_size; // @[SimTop.scala 23:17]
  assign dcache_io_dmem_data_strb = core_io_dmem_data_strb; // @[SimTop.scala 23:17]
  assign dcache_io_dmem_data_write = core_io_dmem_data_write; // @[SimTop.scala 23:17]
  assign dcache_io_out_data_ready = top_io_dmem_data_ready; // @[SimTop.scala 24:17]
  assign dcache_io_out_data_read = top_io_dmem_data_read; // @[SimTop.scala 24:17]
  assign top_clock = clock;
  assign top_reset = reset;
  assign top_io_out_aw_ready = io_memAXI_0_aw_ready; // @[SimTop.scala 33:18]
  assign top_io_out_w_ready = io_memAXI_0_w_ready; // @[SimTop.scala 34:18]
  assign top_io_out_b_valid = io_memAXI_0_b_valid; // @[SimTop.scala 35:18]
  assign top_io_out_ar_ready = io_memAXI_0_ar_ready; // @[SimTop.scala 36:18]
  assign top_io_out_r_valid = io_memAXI_0_r_valid; // @[SimTop.scala 37:18]
  assign top_io_out_r_bits_data = io_memAXI_0_r_bits_data; // @[SimTop.scala 37:18]
  assign top_io_out_r_bits_last = io_memAXI_0_r_bits_last; // @[SimTop.scala 37:18]
  assign top_io_imem_inst_valid = icache_io_out_inst_valid; // @[SimTop.scala 22:17]
  assign top_io_imem_inst_addr = icache_io_out_inst_addr; // @[SimTop.scala 22:17]
  assign top_io_dmem_data_valid = dcache_io_out_data_valid; // @[SimTop.scala 24:17]
  assign top_io_dmem_data_req = dcache_io_out_data_req; // @[SimTop.scala 24:17]
  assign top_io_dmem_data_addr = dcache_io_out_data_addr; // @[SimTop.scala 24:17]
  assign top_io_dmem_data_strb = dcache_io_out_data_strb; // @[SimTop.scala 24:17]
  assign top_io_dmem_data_write = dcache_io_out_data_write; // @[SimTop.scala 24:17]
endmodule
