module BrPredictor(
  input         clock,
  input         reset,
  input  [31:0] io_pc,
  input         io_is_br,
  input         io_jmp_packet_valid,
  input  [31:0] io_jmp_packet_inst_pc,
  input         io_jmp_packet_jmp,
  input  [31:0] io_jmp_packet_jmp_pc,
  input         io_jmp_packet_mis,
  output        io_pred_br,
  output [31:0] io_pred_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [31:0] _RAND_2187;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [31:0] _RAND_2193;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2202;
  reg [31:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2218;
  reg [31:0] _RAND_2219;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [31:0] _RAND_2241;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2245;
  reg [31:0] _RAND_2246;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [31:0] _RAND_2265;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [31:0] _RAND_2271;
  reg [31:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2281;
  reg [31:0] _RAND_2282;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] npc = io_pc + 32'h4; // @[BrPredictor.scala 39:19]
  reg [5:0] bht_0; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_1; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_2; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_3; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_4; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_5; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_6; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_7; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_8; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_9; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_10; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_11; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_12; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_13; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_14; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_15; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_16; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_17; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_18; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_19; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_20; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_21; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_22; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_23; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_24; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_25; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_26; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_27; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_28; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_29; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_30; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_31; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_32; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_33; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_34; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_35; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_36; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_37; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_38; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_39; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_40; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_41; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_42; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_43; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_44; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_45; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_46; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_47; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_48; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_49; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_50; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_51; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_52; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_53; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_54; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_55; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_56; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_57; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_58; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_59; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_60; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_61; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_62; // @[BrPredictor.scala 50:20]
  reg [5:0] bht_63; // @[BrPredictor.scala 50:20]
  reg [1:0] pht_0_0; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_1; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_2; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_3; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_4; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_5; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_6; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_7; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_8; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_9; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_10; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_11; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_12; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_13; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_14; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_15; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_16; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_17; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_18; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_19; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_20; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_21; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_22; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_23; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_24; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_25; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_26; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_27; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_28; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_29; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_30; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_31; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_32; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_33; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_34; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_35; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_36; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_37; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_38; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_39; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_40; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_41; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_42; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_43; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_44; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_45; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_46; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_47; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_48; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_49; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_50; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_51; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_52; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_53; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_54; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_55; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_56; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_57; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_58; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_59; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_60; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_61; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_62; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_63; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_64; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_65; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_66; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_67; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_68; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_69; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_70; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_71; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_72; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_73; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_74; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_75; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_76; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_77; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_78; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_79; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_80; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_81; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_82; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_83; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_84; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_85; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_86; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_87; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_88; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_89; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_90; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_91; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_92; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_93; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_94; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_95; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_96; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_97; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_98; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_99; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_100; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_101; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_102; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_103; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_104; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_105; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_106; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_107; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_108; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_109; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_110; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_111; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_112; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_113; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_114; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_115; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_116; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_117; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_118; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_119; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_120; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_121; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_122; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_123; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_124; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_125; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_126; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_127; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_128; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_129; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_130; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_131; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_132; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_133; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_134; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_135; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_136; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_137; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_138; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_139; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_140; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_141; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_142; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_143; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_144; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_145; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_146; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_147; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_148; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_149; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_150; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_151; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_152; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_153; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_154; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_155; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_156; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_157; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_158; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_159; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_160; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_161; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_162; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_163; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_164; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_165; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_166; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_167; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_168; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_169; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_170; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_171; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_172; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_173; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_174; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_175; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_176; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_177; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_178; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_179; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_180; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_181; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_182; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_183; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_184; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_185; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_186; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_187; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_188; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_189; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_190; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_191; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_192; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_193; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_194; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_195; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_196; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_197; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_198; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_199; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_200; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_201; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_202; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_203; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_204; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_205; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_206; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_207; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_208; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_209; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_210; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_211; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_212; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_213; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_214; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_215; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_216; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_217; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_218; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_219; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_220; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_221; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_222; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_223; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_224; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_225; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_226; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_227; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_228; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_229; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_230; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_231; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_232; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_233; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_234; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_235; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_236; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_237; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_238; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_239; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_240; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_241; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_242; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_243; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_244; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_245; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_246; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_247; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_248; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_249; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_250; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_251; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_252; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_253; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_254; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_0_255; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_0; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_1; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_2; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_3; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_4; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_5; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_6; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_7; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_8; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_9; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_10; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_11; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_12; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_13; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_14; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_15; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_16; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_17; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_18; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_19; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_20; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_21; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_22; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_23; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_24; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_25; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_26; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_27; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_28; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_29; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_30; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_31; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_32; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_33; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_34; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_35; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_36; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_37; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_38; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_39; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_40; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_41; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_42; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_43; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_44; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_45; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_46; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_47; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_48; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_49; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_50; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_51; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_52; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_53; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_54; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_55; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_56; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_57; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_58; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_59; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_60; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_61; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_62; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_63; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_64; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_65; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_66; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_67; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_68; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_69; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_70; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_71; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_72; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_73; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_74; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_75; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_76; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_77; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_78; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_79; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_80; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_81; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_82; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_83; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_84; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_85; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_86; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_87; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_88; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_89; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_90; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_91; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_92; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_93; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_94; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_95; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_96; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_97; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_98; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_99; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_100; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_101; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_102; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_103; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_104; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_105; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_106; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_107; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_108; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_109; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_110; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_111; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_112; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_113; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_114; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_115; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_116; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_117; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_118; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_119; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_120; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_121; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_122; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_123; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_124; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_125; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_126; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_127; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_128; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_129; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_130; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_131; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_132; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_133; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_134; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_135; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_136; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_137; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_138; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_139; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_140; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_141; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_142; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_143; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_144; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_145; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_146; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_147; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_148; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_149; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_150; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_151; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_152; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_153; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_154; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_155; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_156; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_157; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_158; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_159; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_160; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_161; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_162; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_163; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_164; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_165; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_166; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_167; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_168; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_169; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_170; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_171; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_172; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_173; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_174; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_175; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_176; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_177; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_178; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_179; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_180; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_181; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_182; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_183; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_184; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_185; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_186; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_187; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_188; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_189; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_190; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_191; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_192; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_193; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_194; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_195; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_196; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_197; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_198; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_199; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_200; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_201; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_202; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_203; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_204; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_205; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_206; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_207; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_208; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_209; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_210; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_211; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_212; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_213; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_214; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_215; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_216; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_217; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_218; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_219; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_220; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_221; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_222; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_223; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_224; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_225; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_226; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_227; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_228; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_229; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_230; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_231; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_232; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_233; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_234; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_235; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_236; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_237; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_238; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_239; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_240; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_241; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_242; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_243; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_244; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_245; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_246; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_247; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_248; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_249; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_250; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_251; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_252; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_253; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_254; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_1_255; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_0; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_1; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_2; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_3; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_4; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_5; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_6; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_7; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_8; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_9; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_10; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_11; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_12; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_13; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_14; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_15; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_16; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_17; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_18; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_19; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_20; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_21; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_22; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_23; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_24; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_25; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_26; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_27; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_28; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_29; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_30; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_31; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_32; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_33; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_34; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_35; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_36; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_37; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_38; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_39; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_40; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_41; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_42; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_43; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_44; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_45; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_46; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_47; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_48; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_49; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_50; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_51; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_52; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_53; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_54; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_55; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_56; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_57; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_58; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_59; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_60; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_61; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_62; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_63; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_64; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_65; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_66; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_67; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_68; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_69; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_70; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_71; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_72; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_73; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_74; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_75; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_76; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_77; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_78; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_79; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_80; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_81; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_82; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_83; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_84; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_85; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_86; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_87; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_88; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_89; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_90; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_91; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_92; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_93; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_94; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_95; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_96; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_97; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_98; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_99; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_100; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_101; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_102; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_103; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_104; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_105; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_106; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_107; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_108; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_109; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_110; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_111; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_112; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_113; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_114; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_115; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_116; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_117; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_118; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_119; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_120; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_121; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_122; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_123; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_124; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_125; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_126; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_127; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_128; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_129; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_130; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_131; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_132; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_133; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_134; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_135; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_136; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_137; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_138; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_139; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_140; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_141; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_142; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_143; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_144; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_145; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_146; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_147; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_148; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_149; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_150; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_151; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_152; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_153; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_154; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_155; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_156; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_157; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_158; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_159; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_160; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_161; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_162; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_163; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_164; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_165; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_166; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_167; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_168; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_169; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_170; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_171; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_172; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_173; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_174; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_175; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_176; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_177; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_178; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_179; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_180; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_181; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_182; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_183; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_184; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_185; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_186; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_187; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_188; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_189; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_190; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_191; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_192; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_193; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_194; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_195; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_196; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_197; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_198; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_199; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_200; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_201; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_202; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_203; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_204; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_205; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_206; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_207; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_208; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_209; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_210; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_211; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_212; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_213; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_214; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_215; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_216; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_217; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_218; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_219; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_220; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_221; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_222; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_223; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_224; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_225; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_226; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_227; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_228; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_229; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_230; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_231; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_232; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_233; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_234; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_235; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_236; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_237; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_238; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_239; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_240; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_241; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_242; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_243; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_244; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_245; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_246; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_247; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_248; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_249; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_250; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_251; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_252; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_253; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_254; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_2_255; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_0; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_1; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_2; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_3; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_4; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_5; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_6; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_7; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_8; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_9; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_10; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_11; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_12; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_13; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_14; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_15; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_16; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_17; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_18; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_19; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_20; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_21; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_22; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_23; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_24; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_25; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_26; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_27; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_28; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_29; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_30; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_31; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_32; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_33; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_34; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_35; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_36; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_37; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_38; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_39; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_40; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_41; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_42; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_43; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_44; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_45; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_46; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_47; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_48; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_49; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_50; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_51; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_52; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_53; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_54; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_55; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_56; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_57; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_58; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_59; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_60; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_61; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_62; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_63; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_64; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_65; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_66; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_67; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_68; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_69; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_70; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_71; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_72; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_73; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_74; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_75; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_76; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_77; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_78; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_79; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_80; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_81; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_82; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_83; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_84; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_85; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_86; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_87; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_88; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_89; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_90; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_91; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_92; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_93; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_94; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_95; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_96; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_97; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_98; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_99; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_100; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_101; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_102; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_103; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_104; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_105; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_106; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_107; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_108; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_109; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_110; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_111; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_112; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_113; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_114; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_115; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_116; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_117; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_118; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_119; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_120; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_121; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_122; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_123; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_124; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_125; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_126; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_127; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_128; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_129; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_130; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_131; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_132; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_133; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_134; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_135; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_136; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_137; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_138; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_139; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_140; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_141; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_142; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_143; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_144; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_145; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_146; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_147; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_148; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_149; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_150; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_151; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_152; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_153; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_154; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_155; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_156; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_157; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_158; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_159; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_160; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_161; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_162; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_163; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_164; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_165; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_166; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_167; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_168; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_169; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_170; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_171; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_172; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_173; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_174; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_175; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_176; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_177; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_178; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_179; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_180; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_181; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_182; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_183; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_184; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_185; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_186; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_187; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_188; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_189; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_190; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_191; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_192; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_193; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_194; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_195; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_196; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_197; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_198; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_199; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_200; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_201; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_202; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_203; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_204; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_205; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_206; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_207; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_208; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_209; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_210; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_211; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_212; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_213; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_214; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_215; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_216; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_217; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_218; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_219; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_220; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_221; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_222; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_223; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_224; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_225; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_226; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_227; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_228; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_229; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_230; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_231; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_232; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_233; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_234; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_235; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_236; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_237; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_238; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_239; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_240; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_241; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_242; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_243; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_244; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_245; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_246; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_247; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_248; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_249; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_250; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_251; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_252; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_253; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_254; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_3_255; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_0; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_1; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_2; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_3; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_4; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_5; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_6; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_7; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_8; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_9; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_10; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_11; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_12; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_13; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_14; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_15; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_16; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_17; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_18; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_19; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_20; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_21; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_22; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_23; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_24; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_25; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_26; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_27; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_28; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_29; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_30; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_31; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_32; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_33; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_34; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_35; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_36; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_37; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_38; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_39; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_40; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_41; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_42; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_43; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_44; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_45; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_46; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_47; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_48; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_49; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_50; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_51; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_52; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_53; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_54; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_55; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_56; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_57; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_58; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_59; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_60; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_61; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_62; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_63; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_64; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_65; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_66; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_67; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_68; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_69; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_70; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_71; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_72; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_73; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_74; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_75; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_76; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_77; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_78; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_79; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_80; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_81; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_82; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_83; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_84; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_85; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_86; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_87; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_88; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_89; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_90; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_91; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_92; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_93; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_94; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_95; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_96; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_97; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_98; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_99; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_100; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_101; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_102; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_103; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_104; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_105; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_106; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_107; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_108; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_109; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_110; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_111; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_112; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_113; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_114; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_115; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_116; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_117; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_118; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_119; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_120; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_121; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_122; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_123; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_124; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_125; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_126; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_127; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_128; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_129; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_130; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_131; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_132; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_133; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_134; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_135; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_136; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_137; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_138; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_139; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_140; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_141; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_142; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_143; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_144; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_145; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_146; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_147; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_148; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_149; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_150; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_151; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_152; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_153; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_154; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_155; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_156; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_157; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_158; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_159; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_160; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_161; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_162; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_163; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_164; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_165; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_166; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_167; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_168; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_169; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_170; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_171; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_172; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_173; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_174; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_175; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_176; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_177; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_178; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_179; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_180; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_181; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_182; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_183; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_184; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_185; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_186; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_187; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_188; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_189; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_190; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_191; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_192; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_193; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_194; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_195; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_196; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_197; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_198; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_199; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_200; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_201; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_202; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_203; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_204; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_205; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_206; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_207; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_208; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_209; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_210; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_211; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_212; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_213; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_214; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_215; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_216; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_217; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_218; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_219; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_220; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_221; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_222; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_223; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_224; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_225; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_226; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_227; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_228; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_229; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_230; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_231; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_232; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_233; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_234; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_235; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_236; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_237; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_238; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_239; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_240; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_241; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_242; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_243; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_244; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_245; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_246; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_247; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_248; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_249; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_250; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_251; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_252; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_253; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_254; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_4_255; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_0; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_1; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_2; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_3; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_4; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_5; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_6; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_7; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_8; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_9; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_10; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_11; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_12; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_13; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_14; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_15; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_16; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_17; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_18; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_19; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_20; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_21; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_22; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_23; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_24; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_25; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_26; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_27; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_28; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_29; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_30; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_31; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_32; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_33; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_34; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_35; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_36; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_37; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_38; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_39; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_40; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_41; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_42; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_43; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_44; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_45; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_46; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_47; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_48; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_49; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_50; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_51; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_52; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_53; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_54; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_55; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_56; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_57; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_58; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_59; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_60; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_61; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_62; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_63; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_64; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_65; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_66; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_67; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_68; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_69; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_70; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_71; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_72; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_73; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_74; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_75; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_76; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_77; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_78; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_79; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_80; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_81; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_82; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_83; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_84; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_85; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_86; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_87; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_88; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_89; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_90; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_91; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_92; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_93; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_94; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_95; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_96; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_97; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_98; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_99; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_100; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_101; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_102; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_103; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_104; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_105; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_106; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_107; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_108; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_109; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_110; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_111; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_112; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_113; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_114; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_115; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_116; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_117; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_118; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_119; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_120; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_121; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_122; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_123; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_124; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_125; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_126; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_127; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_128; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_129; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_130; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_131; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_132; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_133; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_134; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_135; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_136; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_137; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_138; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_139; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_140; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_141; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_142; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_143; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_144; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_145; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_146; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_147; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_148; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_149; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_150; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_151; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_152; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_153; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_154; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_155; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_156; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_157; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_158; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_159; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_160; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_161; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_162; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_163; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_164; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_165; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_166; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_167; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_168; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_169; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_170; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_171; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_172; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_173; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_174; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_175; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_176; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_177; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_178; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_179; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_180; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_181; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_182; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_183; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_184; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_185; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_186; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_187; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_188; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_189; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_190; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_191; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_192; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_193; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_194; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_195; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_196; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_197; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_198; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_199; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_200; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_201; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_202; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_203; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_204; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_205; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_206; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_207; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_208; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_209; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_210; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_211; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_212; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_213; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_214; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_215; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_216; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_217; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_218; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_219; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_220; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_221; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_222; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_223; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_224; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_225; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_226; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_227; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_228; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_229; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_230; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_231; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_232; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_233; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_234; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_235; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_236; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_237; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_238; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_239; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_240; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_241; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_242; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_243; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_244; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_245; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_246; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_247; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_248; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_249; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_250; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_251; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_252; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_253; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_254; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_5_255; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_0; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_1; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_2; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_3; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_4; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_5; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_6; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_7; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_8; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_9; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_10; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_11; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_12; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_13; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_14; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_15; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_16; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_17; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_18; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_19; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_20; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_21; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_22; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_23; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_24; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_25; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_26; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_27; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_28; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_29; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_30; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_31; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_32; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_33; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_34; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_35; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_36; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_37; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_38; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_39; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_40; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_41; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_42; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_43; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_44; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_45; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_46; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_47; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_48; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_49; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_50; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_51; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_52; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_53; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_54; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_55; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_56; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_57; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_58; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_59; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_60; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_61; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_62; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_63; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_64; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_65; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_66; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_67; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_68; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_69; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_70; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_71; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_72; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_73; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_74; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_75; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_76; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_77; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_78; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_79; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_80; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_81; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_82; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_83; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_84; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_85; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_86; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_87; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_88; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_89; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_90; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_91; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_92; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_93; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_94; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_95; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_96; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_97; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_98; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_99; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_100; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_101; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_102; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_103; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_104; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_105; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_106; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_107; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_108; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_109; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_110; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_111; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_112; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_113; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_114; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_115; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_116; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_117; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_118; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_119; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_120; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_121; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_122; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_123; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_124; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_125; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_126; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_127; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_128; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_129; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_130; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_131; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_132; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_133; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_134; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_135; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_136; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_137; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_138; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_139; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_140; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_141; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_142; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_143; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_144; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_145; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_146; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_147; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_148; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_149; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_150; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_151; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_152; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_153; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_154; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_155; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_156; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_157; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_158; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_159; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_160; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_161; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_162; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_163; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_164; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_165; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_166; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_167; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_168; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_169; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_170; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_171; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_172; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_173; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_174; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_175; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_176; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_177; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_178; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_179; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_180; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_181; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_182; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_183; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_184; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_185; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_186; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_187; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_188; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_189; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_190; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_191; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_192; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_193; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_194; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_195; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_196; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_197; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_198; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_199; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_200; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_201; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_202; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_203; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_204; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_205; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_206; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_207; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_208; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_209; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_210; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_211; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_212; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_213; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_214; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_215; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_216; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_217; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_218; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_219; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_220; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_221; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_222; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_223; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_224; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_225; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_226; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_227; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_228; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_229; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_230; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_231; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_232; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_233; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_234; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_235; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_236; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_237; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_238; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_239; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_240; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_241; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_242; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_243; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_244; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_245; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_246; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_247; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_248; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_249; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_250; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_251; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_252; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_253; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_254; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_6_255; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_0; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_1; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_2; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_3; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_4; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_5; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_6; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_7; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_8; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_9; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_10; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_11; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_12; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_13; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_14; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_15; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_16; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_17; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_18; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_19; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_20; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_21; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_22; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_23; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_24; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_25; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_26; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_27; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_28; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_29; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_30; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_31; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_32; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_33; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_34; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_35; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_36; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_37; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_38; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_39; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_40; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_41; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_42; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_43; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_44; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_45; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_46; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_47; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_48; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_49; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_50; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_51; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_52; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_53; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_54; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_55; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_56; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_57; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_58; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_59; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_60; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_61; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_62; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_63; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_64; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_65; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_66; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_67; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_68; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_69; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_70; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_71; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_72; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_73; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_74; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_75; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_76; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_77; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_78; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_79; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_80; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_81; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_82; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_83; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_84; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_85; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_86; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_87; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_88; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_89; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_90; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_91; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_92; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_93; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_94; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_95; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_96; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_97; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_98; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_99; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_100; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_101; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_102; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_103; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_104; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_105; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_106; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_107; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_108; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_109; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_110; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_111; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_112; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_113; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_114; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_115; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_116; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_117; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_118; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_119; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_120; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_121; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_122; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_123; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_124; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_125; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_126; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_127; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_128; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_129; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_130; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_131; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_132; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_133; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_134; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_135; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_136; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_137; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_138; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_139; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_140; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_141; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_142; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_143; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_144; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_145; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_146; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_147; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_148; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_149; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_150; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_151; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_152; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_153; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_154; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_155; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_156; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_157; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_158; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_159; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_160; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_161; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_162; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_163; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_164; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_165; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_166; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_167; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_168; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_169; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_170; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_171; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_172; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_173; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_174; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_175; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_176; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_177; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_178; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_179; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_180; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_181; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_182; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_183; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_184; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_185; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_186; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_187; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_188; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_189; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_190; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_191; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_192; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_193; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_194; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_195; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_196; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_197; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_198; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_199; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_200; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_201; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_202; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_203; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_204; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_205; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_206; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_207; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_208; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_209; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_210; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_211; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_212; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_213; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_214; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_215; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_216; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_217; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_218; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_219; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_220; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_221; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_222; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_223; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_224; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_225; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_226; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_227; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_228; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_229; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_230; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_231; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_232; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_233; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_234; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_235; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_236; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_237; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_238; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_239; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_240; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_241; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_242; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_243; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_244; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_245; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_246; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_247; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_248; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_249; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_250; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_251; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_252; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_253; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_254; // @[BrPredictor.scala 51:20]
  reg [1:0] pht_7_255; // @[BrPredictor.scala 51:20]
  wire [5:0] bht_raddr = io_pc[7:2]; // @[BrPredictor.scala 52:34]
  wire [5:0] _GEN_1 = 6'h1 == bht_raddr ? bht_1 : bht_0; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_2 = 6'h2 == bht_raddr ? bht_2 : _GEN_1; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_3 = 6'h3 == bht_raddr ? bht_3 : _GEN_2; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_4 = 6'h4 == bht_raddr ? bht_4 : _GEN_3; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_5 = 6'h5 == bht_raddr ? bht_5 : _GEN_4; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_6 = 6'h6 == bht_raddr ? bht_6 : _GEN_5; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_7 = 6'h7 == bht_raddr ? bht_7 : _GEN_6; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_8 = 6'h8 == bht_raddr ? bht_8 : _GEN_7; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_9 = 6'h9 == bht_raddr ? bht_9 : _GEN_8; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_10 = 6'ha == bht_raddr ? bht_10 : _GEN_9; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_11 = 6'hb == bht_raddr ? bht_11 : _GEN_10; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_12 = 6'hc == bht_raddr ? bht_12 : _GEN_11; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_13 = 6'hd == bht_raddr ? bht_13 : _GEN_12; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_14 = 6'he == bht_raddr ? bht_14 : _GEN_13; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_15 = 6'hf == bht_raddr ? bht_15 : _GEN_14; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_16 = 6'h10 == bht_raddr ? bht_16 : _GEN_15; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_17 = 6'h11 == bht_raddr ? bht_17 : _GEN_16; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_18 = 6'h12 == bht_raddr ? bht_18 : _GEN_17; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_19 = 6'h13 == bht_raddr ? bht_19 : _GEN_18; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_20 = 6'h14 == bht_raddr ? bht_20 : _GEN_19; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_21 = 6'h15 == bht_raddr ? bht_21 : _GEN_20; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_22 = 6'h16 == bht_raddr ? bht_22 : _GEN_21; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_23 = 6'h17 == bht_raddr ? bht_23 : _GEN_22; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_24 = 6'h18 == bht_raddr ? bht_24 : _GEN_23; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_25 = 6'h19 == bht_raddr ? bht_25 : _GEN_24; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_26 = 6'h1a == bht_raddr ? bht_26 : _GEN_25; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_27 = 6'h1b == bht_raddr ? bht_27 : _GEN_26; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_28 = 6'h1c == bht_raddr ? bht_28 : _GEN_27; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_29 = 6'h1d == bht_raddr ? bht_29 : _GEN_28; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_30 = 6'h1e == bht_raddr ? bht_30 : _GEN_29; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_31 = 6'h1f == bht_raddr ? bht_31 : _GEN_30; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_32 = 6'h20 == bht_raddr ? bht_32 : _GEN_31; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_33 = 6'h21 == bht_raddr ? bht_33 : _GEN_32; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_34 = 6'h22 == bht_raddr ? bht_34 : _GEN_33; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_35 = 6'h23 == bht_raddr ? bht_35 : _GEN_34; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_36 = 6'h24 == bht_raddr ? bht_36 : _GEN_35; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_37 = 6'h25 == bht_raddr ? bht_37 : _GEN_36; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_38 = 6'h26 == bht_raddr ? bht_38 : _GEN_37; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_39 = 6'h27 == bht_raddr ? bht_39 : _GEN_38; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_40 = 6'h28 == bht_raddr ? bht_40 : _GEN_39; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_41 = 6'h29 == bht_raddr ? bht_41 : _GEN_40; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_42 = 6'h2a == bht_raddr ? bht_42 : _GEN_41; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_43 = 6'h2b == bht_raddr ? bht_43 : _GEN_42; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_44 = 6'h2c == bht_raddr ? bht_44 : _GEN_43; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_45 = 6'h2d == bht_raddr ? bht_45 : _GEN_44; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_46 = 6'h2e == bht_raddr ? bht_46 : _GEN_45; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_47 = 6'h2f == bht_raddr ? bht_47 : _GEN_46; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_48 = 6'h30 == bht_raddr ? bht_48 : _GEN_47; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_49 = 6'h31 == bht_raddr ? bht_49 : _GEN_48; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_50 = 6'h32 == bht_raddr ? bht_50 : _GEN_49; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_51 = 6'h33 == bht_raddr ? bht_51 : _GEN_50; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_52 = 6'h34 == bht_raddr ? bht_52 : _GEN_51; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_53 = 6'h35 == bht_raddr ? bht_53 : _GEN_52; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_54 = 6'h36 == bht_raddr ? bht_54 : _GEN_53; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_55 = 6'h37 == bht_raddr ? bht_55 : _GEN_54; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_56 = 6'h38 == bht_raddr ? bht_56 : _GEN_55; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_57 = 6'h39 == bht_raddr ? bht_57 : _GEN_56; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_58 = 6'h3a == bht_raddr ? bht_58 : _GEN_57; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_59 = 6'h3b == bht_raddr ? bht_59 : _GEN_58; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_60 = 6'h3c == bht_raddr ? bht_60 : _GEN_59; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_61 = 6'h3d == bht_raddr ? bht_61 : _GEN_60; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_62 = 6'h3e == bht_raddr ? bht_62 : _GEN_61; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] _GEN_63 = 6'h3f == bht_raddr ? bht_63 : _GEN_62; // @[BrPredictor.scala 53:58 BrPredictor.scala 53:58]
  wire [5:0] pht_raddr = _GEN_63 ^ bht_raddr; // @[BrPredictor.scala 53:58]
  wire [2:0] pht_rindex = io_pc[10:8]; // @[BrPredictor.scala 54:35]
  wire [1:0] _GEN_65 = 3'h0 == pht_rindex & 6'h1 == pht_raddr ? pht_0_1 : pht_0_0; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_66 = 3'h0 == pht_rindex & 6'h2 == pht_raddr ? pht_0_2 : _GEN_65; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_67 = 3'h0 == pht_rindex & 6'h3 == pht_raddr ? pht_0_3 : _GEN_66; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_68 = 3'h0 == pht_rindex & 6'h4 == pht_raddr ? pht_0_4 : _GEN_67; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_69 = 3'h0 == pht_rindex & 6'h5 == pht_raddr ? pht_0_5 : _GEN_68; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_70 = 3'h0 == pht_rindex & 6'h6 == pht_raddr ? pht_0_6 : _GEN_69; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_71 = 3'h0 == pht_rindex & 6'h7 == pht_raddr ? pht_0_7 : _GEN_70; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_72 = 3'h0 == pht_rindex & 6'h8 == pht_raddr ? pht_0_8 : _GEN_71; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_73 = 3'h0 == pht_rindex & 6'h9 == pht_raddr ? pht_0_9 : _GEN_72; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_74 = 3'h0 == pht_rindex & 6'ha == pht_raddr ? pht_0_10 : _GEN_73; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_75 = 3'h0 == pht_rindex & 6'hb == pht_raddr ? pht_0_11 : _GEN_74; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_76 = 3'h0 == pht_rindex & 6'hc == pht_raddr ? pht_0_12 : _GEN_75; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_77 = 3'h0 == pht_rindex & 6'hd == pht_raddr ? pht_0_13 : _GEN_76; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_78 = 3'h0 == pht_rindex & 6'he == pht_raddr ? pht_0_14 : _GEN_77; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_79 = 3'h0 == pht_rindex & 6'hf == pht_raddr ? pht_0_15 : _GEN_78; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_80 = 3'h0 == pht_rindex & 6'h10 == pht_raddr ? pht_0_16 : _GEN_79; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_81 = 3'h0 == pht_rindex & 6'h11 == pht_raddr ? pht_0_17 : _GEN_80; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_82 = 3'h0 == pht_rindex & 6'h12 == pht_raddr ? pht_0_18 : _GEN_81; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_83 = 3'h0 == pht_rindex & 6'h13 == pht_raddr ? pht_0_19 : _GEN_82; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_84 = 3'h0 == pht_rindex & 6'h14 == pht_raddr ? pht_0_20 : _GEN_83; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_85 = 3'h0 == pht_rindex & 6'h15 == pht_raddr ? pht_0_21 : _GEN_84; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_86 = 3'h0 == pht_rindex & 6'h16 == pht_raddr ? pht_0_22 : _GEN_85; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_87 = 3'h0 == pht_rindex & 6'h17 == pht_raddr ? pht_0_23 : _GEN_86; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_88 = 3'h0 == pht_rindex & 6'h18 == pht_raddr ? pht_0_24 : _GEN_87; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_89 = 3'h0 == pht_rindex & 6'h19 == pht_raddr ? pht_0_25 : _GEN_88; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_90 = 3'h0 == pht_rindex & 6'h1a == pht_raddr ? pht_0_26 : _GEN_89; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_91 = 3'h0 == pht_rindex & 6'h1b == pht_raddr ? pht_0_27 : _GEN_90; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_92 = 3'h0 == pht_rindex & 6'h1c == pht_raddr ? pht_0_28 : _GEN_91; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_93 = 3'h0 == pht_rindex & 6'h1d == pht_raddr ? pht_0_29 : _GEN_92; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_94 = 3'h0 == pht_rindex & 6'h1e == pht_raddr ? pht_0_30 : _GEN_93; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_95 = 3'h0 == pht_rindex & 6'h1f == pht_raddr ? pht_0_31 : _GEN_94; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_96 = 3'h0 == pht_rindex & 6'h20 == pht_raddr ? pht_0_32 : _GEN_95; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_97 = 3'h0 == pht_rindex & 6'h21 == pht_raddr ? pht_0_33 : _GEN_96; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_98 = 3'h0 == pht_rindex & 6'h22 == pht_raddr ? pht_0_34 : _GEN_97; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_99 = 3'h0 == pht_rindex & 6'h23 == pht_raddr ? pht_0_35 : _GEN_98; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_100 = 3'h0 == pht_rindex & 6'h24 == pht_raddr ? pht_0_36 : _GEN_99; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_101 = 3'h0 == pht_rindex & 6'h25 == pht_raddr ? pht_0_37 : _GEN_100; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_102 = 3'h0 == pht_rindex & 6'h26 == pht_raddr ? pht_0_38 : _GEN_101; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_103 = 3'h0 == pht_rindex & 6'h27 == pht_raddr ? pht_0_39 : _GEN_102; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_104 = 3'h0 == pht_rindex & 6'h28 == pht_raddr ? pht_0_40 : _GEN_103; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_105 = 3'h0 == pht_rindex & 6'h29 == pht_raddr ? pht_0_41 : _GEN_104; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_106 = 3'h0 == pht_rindex & 6'h2a == pht_raddr ? pht_0_42 : _GEN_105; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_107 = 3'h0 == pht_rindex & 6'h2b == pht_raddr ? pht_0_43 : _GEN_106; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_108 = 3'h0 == pht_rindex & 6'h2c == pht_raddr ? pht_0_44 : _GEN_107; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_109 = 3'h0 == pht_rindex & 6'h2d == pht_raddr ? pht_0_45 : _GEN_108; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_110 = 3'h0 == pht_rindex & 6'h2e == pht_raddr ? pht_0_46 : _GEN_109; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_111 = 3'h0 == pht_rindex & 6'h2f == pht_raddr ? pht_0_47 : _GEN_110; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_112 = 3'h0 == pht_rindex & 6'h30 == pht_raddr ? pht_0_48 : _GEN_111; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_113 = 3'h0 == pht_rindex & 6'h31 == pht_raddr ? pht_0_49 : _GEN_112; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_114 = 3'h0 == pht_rindex & 6'h32 == pht_raddr ? pht_0_50 : _GEN_113; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_115 = 3'h0 == pht_rindex & 6'h33 == pht_raddr ? pht_0_51 : _GEN_114; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_116 = 3'h0 == pht_rindex & 6'h34 == pht_raddr ? pht_0_52 : _GEN_115; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_117 = 3'h0 == pht_rindex & 6'h35 == pht_raddr ? pht_0_53 : _GEN_116; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_118 = 3'h0 == pht_rindex & 6'h36 == pht_raddr ? pht_0_54 : _GEN_117; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_119 = 3'h0 == pht_rindex & 6'h37 == pht_raddr ? pht_0_55 : _GEN_118; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_120 = 3'h0 == pht_rindex & 6'h38 == pht_raddr ? pht_0_56 : _GEN_119; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_121 = 3'h0 == pht_rindex & 6'h39 == pht_raddr ? pht_0_57 : _GEN_120; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_122 = 3'h0 == pht_rindex & 6'h3a == pht_raddr ? pht_0_58 : _GEN_121; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_123 = 3'h0 == pht_rindex & 6'h3b == pht_raddr ? pht_0_59 : _GEN_122; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_124 = 3'h0 == pht_rindex & 6'h3c == pht_raddr ? pht_0_60 : _GEN_123; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_125 = 3'h0 == pht_rindex & 6'h3d == pht_raddr ? pht_0_61 : _GEN_124; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_126 = 3'h0 == pht_rindex & 6'h3e == pht_raddr ? pht_0_62 : _GEN_125; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_127 = 3'h0 == pht_rindex & 6'h3f == pht_raddr ? pht_0_63 : _GEN_126; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [6:0] _GEN_9154 = {{1'd0}, pht_raddr}; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_128 = 3'h0 == pht_rindex & 7'h40 == _GEN_9154 ? pht_0_64 : _GEN_127; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_129 = 3'h0 == pht_rindex & 7'h41 == _GEN_9154 ? pht_0_65 : _GEN_128; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_130 = 3'h0 == pht_rindex & 7'h42 == _GEN_9154 ? pht_0_66 : _GEN_129; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_131 = 3'h0 == pht_rindex & 7'h43 == _GEN_9154 ? pht_0_67 : _GEN_130; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_132 = 3'h0 == pht_rindex & 7'h44 == _GEN_9154 ? pht_0_68 : _GEN_131; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_133 = 3'h0 == pht_rindex & 7'h45 == _GEN_9154 ? pht_0_69 : _GEN_132; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_134 = 3'h0 == pht_rindex & 7'h46 == _GEN_9154 ? pht_0_70 : _GEN_133; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_135 = 3'h0 == pht_rindex & 7'h47 == _GEN_9154 ? pht_0_71 : _GEN_134; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_136 = 3'h0 == pht_rindex & 7'h48 == _GEN_9154 ? pht_0_72 : _GEN_135; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_137 = 3'h0 == pht_rindex & 7'h49 == _GEN_9154 ? pht_0_73 : _GEN_136; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_138 = 3'h0 == pht_rindex & 7'h4a == _GEN_9154 ? pht_0_74 : _GEN_137; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_139 = 3'h0 == pht_rindex & 7'h4b == _GEN_9154 ? pht_0_75 : _GEN_138; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_140 = 3'h0 == pht_rindex & 7'h4c == _GEN_9154 ? pht_0_76 : _GEN_139; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_141 = 3'h0 == pht_rindex & 7'h4d == _GEN_9154 ? pht_0_77 : _GEN_140; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_142 = 3'h0 == pht_rindex & 7'h4e == _GEN_9154 ? pht_0_78 : _GEN_141; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_143 = 3'h0 == pht_rindex & 7'h4f == _GEN_9154 ? pht_0_79 : _GEN_142; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_144 = 3'h0 == pht_rindex & 7'h50 == _GEN_9154 ? pht_0_80 : _GEN_143; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_145 = 3'h0 == pht_rindex & 7'h51 == _GEN_9154 ? pht_0_81 : _GEN_144; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_146 = 3'h0 == pht_rindex & 7'h52 == _GEN_9154 ? pht_0_82 : _GEN_145; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_147 = 3'h0 == pht_rindex & 7'h53 == _GEN_9154 ? pht_0_83 : _GEN_146; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_148 = 3'h0 == pht_rindex & 7'h54 == _GEN_9154 ? pht_0_84 : _GEN_147; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_149 = 3'h0 == pht_rindex & 7'h55 == _GEN_9154 ? pht_0_85 : _GEN_148; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_150 = 3'h0 == pht_rindex & 7'h56 == _GEN_9154 ? pht_0_86 : _GEN_149; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_151 = 3'h0 == pht_rindex & 7'h57 == _GEN_9154 ? pht_0_87 : _GEN_150; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_152 = 3'h0 == pht_rindex & 7'h58 == _GEN_9154 ? pht_0_88 : _GEN_151; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_153 = 3'h0 == pht_rindex & 7'h59 == _GEN_9154 ? pht_0_89 : _GEN_152; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_154 = 3'h0 == pht_rindex & 7'h5a == _GEN_9154 ? pht_0_90 : _GEN_153; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_155 = 3'h0 == pht_rindex & 7'h5b == _GEN_9154 ? pht_0_91 : _GEN_154; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_156 = 3'h0 == pht_rindex & 7'h5c == _GEN_9154 ? pht_0_92 : _GEN_155; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_157 = 3'h0 == pht_rindex & 7'h5d == _GEN_9154 ? pht_0_93 : _GEN_156; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_158 = 3'h0 == pht_rindex & 7'h5e == _GEN_9154 ? pht_0_94 : _GEN_157; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_159 = 3'h0 == pht_rindex & 7'h5f == _GEN_9154 ? pht_0_95 : _GEN_158; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_160 = 3'h0 == pht_rindex & 7'h60 == _GEN_9154 ? pht_0_96 : _GEN_159; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_161 = 3'h0 == pht_rindex & 7'h61 == _GEN_9154 ? pht_0_97 : _GEN_160; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_162 = 3'h0 == pht_rindex & 7'h62 == _GEN_9154 ? pht_0_98 : _GEN_161; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_163 = 3'h0 == pht_rindex & 7'h63 == _GEN_9154 ? pht_0_99 : _GEN_162; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_164 = 3'h0 == pht_rindex & 7'h64 == _GEN_9154 ? pht_0_100 : _GEN_163; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_165 = 3'h0 == pht_rindex & 7'h65 == _GEN_9154 ? pht_0_101 : _GEN_164; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_166 = 3'h0 == pht_rindex & 7'h66 == _GEN_9154 ? pht_0_102 : _GEN_165; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_167 = 3'h0 == pht_rindex & 7'h67 == _GEN_9154 ? pht_0_103 : _GEN_166; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_168 = 3'h0 == pht_rindex & 7'h68 == _GEN_9154 ? pht_0_104 : _GEN_167; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_169 = 3'h0 == pht_rindex & 7'h69 == _GEN_9154 ? pht_0_105 : _GEN_168; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_170 = 3'h0 == pht_rindex & 7'h6a == _GEN_9154 ? pht_0_106 : _GEN_169; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_171 = 3'h0 == pht_rindex & 7'h6b == _GEN_9154 ? pht_0_107 : _GEN_170; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_172 = 3'h0 == pht_rindex & 7'h6c == _GEN_9154 ? pht_0_108 : _GEN_171; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_173 = 3'h0 == pht_rindex & 7'h6d == _GEN_9154 ? pht_0_109 : _GEN_172; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_174 = 3'h0 == pht_rindex & 7'h6e == _GEN_9154 ? pht_0_110 : _GEN_173; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_175 = 3'h0 == pht_rindex & 7'h6f == _GEN_9154 ? pht_0_111 : _GEN_174; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_176 = 3'h0 == pht_rindex & 7'h70 == _GEN_9154 ? pht_0_112 : _GEN_175; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_177 = 3'h0 == pht_rindex & 7'h71 == _GEN_9154 ? pht_0_113 : _GEN_176; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_178 = 3'h0 == pht_rindex & 7'h72 == _GEN_9154 ? pht_0_114 : _GEN_177; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_179 = 3'h0 == pht_rindex & 7'h73 == _GEN_9154 ? pht_0_115 : _GEN_178; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_180 = 3'h0 == pht_rindex & 7'h74 == _GEN_9154 ? pht_0_116 : _GEN_179; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_181 = 3'h0 == pht_rindex & 7'h75 == _GEN_9154 ? pht_0_117 : _GEN_180; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_182 = 3'h0 == pht_rindex & 7'h76 == _GEN_9154 ? pht_0_118 : _GEN_181; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_183 = 3'h0 == pht_rindex & 7'h77 == _GEN_9154 ? pht_0_119 : _GEN_182; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_184 = 3'h0 == pht_rindex & 7'h78 == _GEN_9154 ? pht_0_120 : _GEN_183; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_185 = 3'h0 == pht_rindex & 7'h79 == _GEN_9154 ? pht_0_121 : _GEN_184; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_186 = 3'h0 == pht_rindex & 7'h7a == _GEN_9154 ? pht_0_122 : _GEN_185; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_187 = 3'h0 == pht_rindex & 7'h7b == _GEN_9154 ? pht_0_123 : _GEN_186; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_188 = 3'h0 == pht_rindex & 7'h7c == _GEN_9154 ? pht_0_124 : _GEN_187; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_189 = 3'h0 == pht_rindex & 7'h7d == _GEN_9154 ? pht_0_125 : _GEN_188; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_190 = 3'h0 == pht_rindex & 7'h7e == _GEN_9154 ? pht_0_126 : _GEN_189; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_191 = 3'h0 == pht_rindex & 7'h7f == _GEN_9154 ? pht_0_127 : _GEN_190; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [7:0] _GEN_9346 = {{2'd0}, pht_raddr}; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_192 = 3'h0 == pht_rindex & 8'h80 == _GEN_9346 ? pht_0_128 : _GEN_191; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_193 = 3'h0 == pht_rindex & 8'h81 == _GEN_9346 ? pht_0_129 : _GEN_192; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_194 = 3'h0 == pht_rindex & 8'h82 == _GEN_9346 ? pht_0_130 : _GEN_193; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_195 = 3'h0 == pht_rindex & 8'h83 == _GEN_9346 ? pht_0_131 : _GEN_194; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_196 = 3'h0 == pht_rindex & 8'h84 == _GEN_9346 ? pht_0_132 : _GEN_195; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_197 = 3'h0 == pht_rindex & 8'h85 == _GEN_9346 ? pht_0_133 : _GEN_196; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_198 = 3'h0 == pht_rindex & 8'h86 == _GEN_9346 ? pht_0_134 : _GEN_197; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_199 = 3'h0 == pht_rindex & 8'h87 == _GEN_9346 ? pht_0_135 : _GEN_198; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_200 = 3'h0 == pht_rindex & 8'h88 == _GEN_9346 ? pht_0_136 : _GEN_199; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_201 = 3'h0 == pht_rindex & 8'h89 == _GEN_9346 ? pht_0_137 : _GEN_200; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_202 = 3'h0 == pht_rindex & 8'h8a == _GEN_9346 ? pht_0_138 : _GEN_201; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_203 = 3'h0 == pht_rindex & 8'h8b == _GEN_9346 ? pht_0_139 : _GEN_202; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_204 = 3'h0 == pht_rindex & 8'h8c == _GEN_9346 ? pht_0_140 : _GEN_203; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_205 = 3'h0 == pht_rindex & 8'h8d == _GEN_9346 ? pht_0_141 : _GEN_204; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_206 = 3'h0 == pht_rindex & 8'h8e == _GEN_9346 ? pht_0_142 : _GEN_205; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_207 = 3'h0 == pht_rindex & 8'h8f == _GEN_9346 ? pht_0_143 : _GEN_206; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_208 = 3'h0 == pht_rindex & 8'h90 == _GEN_9346 ? pht_0_144 : _GEN_207; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_209 = 3'h0 == pht_rindex & 8'h91 == _GEN_9346 ? pht_0_145 : _GEN_208; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_210 = 3'h0 == pht_rindex & 8'h92 == _GEN_9346 ? pht_0_146 : _GEN_209; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_211 = 3'h0 == pht_rindex & 8'h93 == _GEN_9346 ? pht_0_147 : _GEN_210; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_212 = 3'h0 == pht_rindex & 8'h94 == _GEN_9346 ? pht_0_148 : _GEN_211; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_213 = 3'h0 == pht_rindex & 8'h95 == _GEN_9346 ? pht_0_149 : _GEN_212; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_214 = 3'h0 == pht_rindex & 8'h96 == _GEN_9346 ? pht_0_150 : _GEN_213; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_215 = 3'h0 == pht_rindex & 8'h97 == _GEN_9346 ? pht_0_151 : _GEN_214; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_216 = 3'h0 == pht_rindex & 8'h98 == _GEN_9346 ? pht_0_152 : _GEN_215; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_217 = 3'h0 == pht_rindex & 8'h99 == _GEN_9346 ? pht_0_153 : _GEN_216; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_218 = 3'h0 == pht_rindex & 8'h9a == _GEN_9346 ? pht_0_154 : _GEN_217; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_219 = 3'h0 == pht_rindex & 8'h9b == _GEN_9346 ? pht_0_155 : _GEN_218; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_220 = 3'h0 == pht_rindex & 8'h9c == _GEN_9346 ? pht_0_156 : _GEN_219; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_221 = 3'h0 == pht_rindex & 8'h9d == _GEN_9346 ? pht_0_157 : _GEN_220; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_222 = 3'h0 == pht_rindex & 8'h9e == _GEN_9346 ? pht_0_158 : _GEN_221; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_223 = 3'h0 == pht_rindex & 8'h9f == _GEN_9346 ? pht_0_159 : _GEN_222; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_224 = 3'h0 == pht_rindex & 8'ha0 == _GEN_9346 ? pht_0_160 : _GEN_223; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_225 = 3'h0 == pht_rindex & 8'ha1 == _GEN_9346 ? pht_0_161 : _GEN_224; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_226 = 3'h0 == pht_rindex & 8'ha2 == _GEN_9346 ? pht_0_162 : _GEN_225; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_227 = 3'h0 == pht_rindex & 8'ha3 == _GEN_9346 ? pht_0_163 : _GEN_226; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_228 = 3'h0 == pht_rindex & 8'ha4 == _GEN_9346 ? pht_0_164 : _GEN_227; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_229 = 3'h0 == pht_rindex & 8'ha5 == _GEN_9346 ? pht_0_165 : _GEN_228; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_230 = 3'h0 == pht_rindex & 8'ha6 == _GEN_9346 ? pht_0_166 : _GEN_229; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_231 = 3'h0 == pht_rindex & 8'ha7 == _GEN_9346 ? pht_0_167 : _GEN_230; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_232 = 3'h0 == pht_rindex & 8'ha8 == _GEN_9346 ? pht_0_168 : _GEN_231; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_233 = 3'h0 == pht_rindex & 8'ha9 == _GEN_9346 ? pht_0_169 : _GEN_232; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_234 = 3'h0 == pht_rindex & 8'haa == _GEN_9346 ? pht_0_170 : _GEN_233; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_235 = 3'h0 == pht_rindex & 8'hab == _GEN_9346 ? pht_0_171 : _GEN_234; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_236 = 3'h0 == pht_rindex & 8'hac == _GEN_9346 ? pht_0_172 : _GEN_235; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_237 = 3'h0 == pht_rindex & 8'had == _GEN_9346 ? pht_0_173 : _GEN_236; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_238 = 3'h0 == pht_rindex & 8'hae == _GEN_9346 ? pht_0_174 : _GEN_237; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_239 = 3'h0 == pht_rindex & 8'haf == _GEN_9346 ? pht_0_175 : _GEN_238; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_240 = 3'h0 == pht_rindex & 8'hb0 == _GEN_9346 ? pht_0_176 : _GEN_239; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_241 = 3'h0 == pht_rindex & 8'hb1 == _GEN_9346 ? pht_0_177 : _GEN_240; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_242 = 3'h0 == pht_rindex & 8'hb2 == _GEN_9346 ? pht_0_178 : _GEN_241; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_243 = 3'h0 == pht_rindex & 8'hb3 == _GEN_9346 ? pht_0_179 : _GEN_242; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_244 = 3'h0 == pht_rindex & 8'hb4 == _GEN_9346 ? pht_0_180 : _GEN_243; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_245 = 3'h0 == pht_rindex & 8'hb5 == _GEN_9346 ? pht_0_181 : _GEN_244; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_246 = 3'h0 == pht_rindex & 8'hb6 == _GEN_9346 ? pht_0_182 : _GEN_245; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_247 = 3'h0 == pht_rindex & 8'hb7 == _GEN_9346 ? pht_0_183 : _GEN_246; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_248 = 3'h0 == pht_rindex & 8'hb8 == _GEN_9346 ? pht_0_184 : _GEN_247; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_249 = 3'h0 == pht_rindex & 8'hb9 == _GEN_9346 ? pht_0_185 : _GEN_248; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_250 = 3'h0 == pht_rindex & 8'hba == _GEN_9346 ? pht_0_186 : _GEN_249; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_251 = 3'h0 == pht_rindex & 8'hbb == _GEN_9346 ? pht_0_187 : _GEN_250; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_252 = 3'h0 == pht_rindex & 8'hbc == _GEN_9346 ? pht_0_188 : _GEN_251; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_253 = 3'h0 == pht_rindex & 8'hbd == _GEN_9346 ? pht_0_189 : _GEN_252; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_254 = 3'h0 == pht_rindex & 8'hbe == _GEN_9346 ? pht_0_190 : _GEN_253; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_255 = 3'h0 == pht_rindex & 8'hbf == _GEN_9346 ? pht_0_191 : _GEN_254; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_256 = 3'h0 == pht_rindex & 8'hc0 == _GEN_9346 ? pht_0_192 : _GEN_255; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_257 = 3'h0 == pht_rindex & 8'hc1 == _GEN_9346 ? pht_0_193 : _GEN_256; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_258 = 3'h0 == pht_rindex & 8'hc2 == _GEN_9346 ? pht_0_194 : _GEN_257; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_259 = 3'h0 == pht_rindex & 8'hc3 == _GEN_9346 ? pht_0_195 : _GEN_258; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_260 = 3'h0 == pht_rindex & 8'hc4 == _GEN_9346 ? pht_0_196 : _GEN_259; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_261 = 3'h0 == pht_rindex & 8'hc5 == _GEN_9346 ? pht_0_197 : _GEN_260; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_262 = 3'h0 == pht_rindex & 8'hc6 == _GEN_9346 ? pht_0_198 : _GEN_261; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_263 = 3'h0 == pht_rindex & 8'hc7 == _GEN_9346 ? pht_0_199 : _GEN_262; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_264 = 3'h0 == pht_rindex & 8'hc8 == _GEN_9346 ? pht_0_200 : _GEN_263; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_265 = 3'h0 == pht_rindex & 8'hc9 == _GEN_9346 ? pht_0_201 : _GEN_264; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_266 = 3'h0 == pht_rindex & 8'hca == _GEN_9346 ? pht_0_202 : _GEN_265; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_267 = 3'h0 == pht_rindex & 8'hcb == _GEN_9346 ? pht_0_203 : _GEN_266; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_268 = 3'h0 == pht_rindex & 8'hcc == _GEN_9346 ? pht_0_204 : _GEN_267; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_269 = 3'h0 == pht_rindex & 8'hcd == _GEN_9346 ? pht_0_205 : _GEN_268; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_270 = 3'h0 == pht_rindex & 8'hce == _GEN_9346 ? pht_0_206 : _GEN_269; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_271 = 3'h0 == pht_rindex & 8'hcf == _GEN_9346 ? pht_0_207 : _GEN_270; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_272 = 3'h0 == pht_rindex & 8'hd0 == _GEN_9346 ? pht_0_208 : _GEN_271; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_273 = 3'h0 == pht_rindex & 8'hd1 == _GEN_9346 ? pht_0_209 : _GEN_272; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_274 = 3'h0 == pht_rindex & 8'hd2 == _GEN_9346 ? pht_0_210 : _GEN_273; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_275 = 3'h0 == pht_rindex & 8'hd3 == _GEN_9346 ? pht_0_211 : _GEN_274; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_276 = 3'h0 == pht_rindex & 8'hd4 == _GEN_9346 ? pht_0_212 : _GEN_275; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_277 = 3'h0 == pht_rindex & 8'hd5 == _GEN_9346 ? pht_0_213 : _GEN_276; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_278 = 3'h0 == pht_rindex & 8'hd6 == _GEN_9346 ? pht_0_214 : _GEN_277; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_279 = 3'h0 == pht_rindex & 8'hd7 == _GEN_9346 ? pht_0_215 : _GEN_278; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_280 = 3'h0 == pht_rindex & 8'hd8 == _GEN_9346 ? pht_0_216 : _GEN_279; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_281 = 3'h0 == pht_rindex & 8'hd9 == _GEN_9346 ? pht_0_217 : _GEN_280; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_282 = 3'h0 == pht_rindex & 8'hda == _GEN_9346 ? pht_0_218 : _GEN_281; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_283 = 3'h0 == pht_rindex & 8'hdb == _GEN_9346 ? pht_0_219 : _GEN_282; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_284 = 3'h0 == pht_rindex & 8'hdc == _GEN_9346 ? pht_0_220 : _GEN_283; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_285 = 3'h0 == pht_rindex & 8'hdd == _GEN_9346 ? pht_0_221 : _GEN_284; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_286 = 3'h0 == pht_rindex & 8'hde == _GEN_9346 ? pht_0_222 : _GEN_285; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_287 = 3'h0 == pht_rindex & 8'hdf == _GEN_9346 ? pht_0_223 : _GEN_286; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_288 = 3'h0 == pht_rindex & 8'he0 == _GEN_9346 ? pht_0_224 : _GEN_287; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_289 = 3'h0 == pht_rindex & 8'he1 == _GEN_9346 ? pht_0_225 : _GEN_288; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_290 = 3'h0 == pht_rindex & 8'he2 == _GEN_9346 ? pht_0_226 : _GEN_289; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_291 = 3'h0 == pht_rindex & 8'he3 == _GEN_9346 ? pht_0_227 : _GEN_290; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_292 = 3'h0 == pht_rindex & 8'he4 == _GEN_9346 ? pht_0_228 : _GEN_291; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_293 = 3'h0 == pht_rindex & 8'he5 == _GEN_9346 ? pht_0_229 : _GEN_292; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_294 = 3'h0 == pht_rindex & 8'he6 == _GEN_9346 ? pht_0_230 : _GEN_293; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_295 = 3'h0 == pht_rindex & 8'he7 == _GEN_9346 ? pht_0_231 : _GEN_294; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_296 = 3'h0 == pht_rindex & 8'he8 == _GEN_9346 ? pht_0_232 : _GEN_295; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_297 = 3'h0 == pht_rindex & 8'he9 == _GEN_9346 ? pht_0_233 : _GEN_296; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_298 = 3'h0 == pht_rindex & 8'hea == _GEN_9346 ? pht_0_234 : _GEN_297; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_299 = 3'h0 == pht_rindex & 8'heb == _GEN_9346 ? pht_0_235 : _GEN_298; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_300 = 3'h0 == pht_rindex & 8'hec == _GEN_9346 ? pht_0_236 : _GEN_299; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_301 = 3'h0 == pht_rindex & 8'hed == _GEN_9346 ? pht_0_237 : _GEN_300; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_302 = 3'h0 == pht_rindex & 8'hee == _GEN_9346 ? pht_0_238 : _GEN_301; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_303 = 3'h0 == pht_rindex & 8'hef == _GEN_9346 ? pht_0_239 : _GEN_302; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_304 = 3'h0 == pht_rindex & 8'hf0 == _GEN_9346 ? pht_0_240 : _GEN_303; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_305 = 3'h0 == pht_rindex & 8'hf1 == _GEN_9346 ? pht_0_241 : _GEN_304; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_306 = 3'h0 == pht_rindex & 8'hf2 == _GEN_9346 ? pht_0_242 : _GEN_305; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_307 = 3'h0 == pht_rindex & 8'hf3 == _GEN_9346 ? pht_0_243 : _GEN_306; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_308 = 3'h0 == pht_rindex & 8'hf4 == _GEN_9346 ? pht_0_244 : _GEN_307; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_309 = 3'h0 == pht_rindex & 8'hf5 == _GEN_9346 ? pht_0_245 : _GEN_308; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_310 = 3'h0 == pht_rindex & 8'hf6 == _GEN_9346 ? pht_0_246 : _GEN_309; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_311 = 3'h0 == pht_rindex & 8'hf7 == _GEN_9346 ? pht_0_247 : _GEN_310; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_312 = 3'h0 == pht_rindex & 8'hf8 == _GEN_9346 ? pht_0_248 : _GEN_311; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_313 = 3'h0 == pht_rindex & 8'hf9 == _GEN_9346 ? pht_0_249 : _GEN_312; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_314 = 3'h0 == pht_rindex & 8'hfa == _GEN_9346 ? pht_0_250 : _GEN_313; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_315 = 3'h0 == pht_rindex & 8'hfb == _GEN_9346 ? pht_0_251 : _GEN_314; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_316 = 3'h0 == pht_rindex & 8'hfc == _GEN_9346 ? pht_0_252 : _GEN_315; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_317 = 3'h0 == pht_rindex & 8'hfd == _GEN_9346 ? pht_0_253 : _GEN_316; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_318 = 3'h0 == pht_rindex & 8'hfe == _GEN_9346 ? pht_0_254 : _GEN_317; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_319 = 3'h0 == pht_rindex & 8'hff == _GEN_9346 ? pht_0_255 : _GEN_318; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_320 = 3'h1 == pht_rindex & 6'h0 == pht_raddr ? pht_1_0 : _GEN_319; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_321 = 3'h1 == pht_rindex & 6'h1 == pht_raddr ? pht_1_1 : _GEN_320; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_322 = 3'h1 == pht_rindex & 6'h2 == pht_raddr ? pht_1_2 : _GEN_321; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_323 = 3'h1 == pht_rindex & 6'h3 == pht_raddr ? pht_1_3 : _GEN_322; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_324 = 3'h1 == pht_rindex & 6'h4 == pht_raddr ? pht_1_4 : _GEN_323; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_325 = 3'h1 == pht_rindex & 6'h5 == pht_raddr ? pht_1_5 : _GEN_324; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_326 = 3'h1 == pht_rindex & 6'h6 == pht_raddr ? pht_1_6 : _GEN_325; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_327 = 3'h1 == pht_rindex & 6'h7 == pht_raddr ? pht_1_7 : _GEN_326; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_328 = 3'h1 == pht_rindex & 6'h8 == pht_raddr ? pht_1_8 : _GEN_327; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_329 = 3'h1 == pht_rindex & 6'h9 == pht_raddr ? pht_1_9 : _GEN_328; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_330 = 3'h1 == pht_rindex & 6'ha == pht_raddr ? pht_1_10 : _GEN_329; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_331 = 3'h1 == pht_rindex & 6'hb == pht_raddr ? pht_1_11 : _GEN_330; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_332 = 3'h1 == pht_rindex & 6'hc == pht_raddr ? pht_1_12 : _GEN_331; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_333 = 3'h1 == pht_rindex & 6'hd == pht_raddr ? pht_1_13 : _GEN_332; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_334 = 3'h1 == pht_rindex & 6'he == pht_raddr ? pht_1_14 : _GEN_333; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_335 = 3'h1 == pht_rindex & 6'hf == pht_raddr ? pht_1_15 : _GEN_334; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_336 = 3'h1 == pht_rindex & 6'h10 == pht_raddr ? pht_1_16 : _GEN_335; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_337 = 3'h1 == pht_rindex & 6'h11 == pht_raddr ? pht_1_17 : _GEN_336; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_338 = 3'h1 == pht_rindex & 6'h12 == pht_raddr ? pht_1_18 : _GEN_337; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_339 = 3'h1 == pht_rindex & 6'h13 == pht_raddr ? pht_1_19 : _GEN_338; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_340 = 3'h1 == pht_rindex & 6'h14 == pht_raddr ? pht_1_20 : _GEN_339; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_341 = 3'h1 == pht_rindex & 6'h15 == pht_raddr ? pht_1_21 : _GEN_340; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_342 = 3'h1 == pht_rindex & 6'h16 == pht_raddr ? pht_1_22 : _GEN_341; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_343 = 3'h1 == pht_rindex & 6'h17 == pht_raddr ? pht_1_23 : _GEN_342; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_344 = 3'h1 == pht_rindex & 6'h18 == pht_raddr ? pht_1_24 : _GEN_343; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_345 = 3'h1 == pht_rindex & 6'h19 == pht_raddr ? pht_1_25 : _GEN_344; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_346 = 3'h1 == pht_rindex & 6'h1a == pht_raddr ? pht_1_26 : _GEN_345; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_347 = 3'h1 == pht_rindex & 6'h1b == pht_raddr ? pht_1_27 : _GEN_346; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_348 = 3'h1 == pht_rindex & 6'h1c == pht_raddr ? pht_1_28 : _GEN_347; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_349 = 3'h1 == pht_rindex & 6'h1d == pht_raddr ? pht_1_29 : _GEN_348; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_350 = 3'h1 == pht_rindex & 6'h1e == pht_raddr ? pht_1_30 : _GEN_349; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_351 = 3'h1 == pht_rindex & 6'h1f == pht_raddr ? pht_1_31 : _GEN_350; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_352 = 3'h1 == pht_rindex & 6'h20 == pht_raddr ? pht_1_32 : _GEN_351; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_353 = 3'h1 == pht_rindex & 6'h21 == pht_raddr ? pht_1_33 : _GEN_352; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_354 = 3'h1 == pht_rindex & 6'h22 == pht_raddr ? pht_1_34 : _GEN_353; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_355 = 3'h1 == pht_rindex & 6'h23 == pht_raddr ? pht_1_35 : _GEN_354; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_356 = 3'h1 == pht_rindex & 6'h24 == pht_raddr ? pht_1_36 : _GEN_355; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_357 = 3'h1 == pht_rindex & 6'h25 == pht_raddr ? pht_1_37 : _GEN_356; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_358 = 3'h1 == pht_rindex & 6'h26 == pht_raddr ? pht_1_38 : _GEN_357; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_359 = 3'h1 == pht_rindex & 6'h27 == pht_raddr ? pht_1_39 : _GEN_358; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_360 = 3'h1 == pht_rindex & 6'h28 == pht_raddr ? pht_1_40 : _GEN_359; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_361 = 3'h1 == pht_rindex & 6'h29 == pht_raddr ? pht_1_41 : _GEN_360; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_362 = 3'h1 == pht_rindex & 6'h2a == pht_raddr ? pht_1_42 : _GEN_361; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_363 = 3'h1 == pht_rindex & 6'h2b == pht_raddr ? pht_1_43 : _GEN_362; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_364 = 3'h1 == pht_rindex & 6'h2c == pht_raddr ? pht_1_44 : _GEN_363; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_365 = 3'h1 == pht_rindex & 6'h2d == pht_raddr ? pht_1_45 : _GEN_364; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_366 = 3'h1 == pht_rindex & 6'h2e == pht_raddr ? pht_1_46 : _GEN_365; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_367 = 3'h1 == pht_rindex & 6'h2f == pht_raddr ? pht_1_47 : _GEN_366; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_368 = 3'h1 == pht_rindex & 6'h30 == pht_raddr ? pht_1_48 : _GEN_367; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_369 = 3'h1 == pht_rindex & 6'h31 == pht_raddr ? pht_1_49 : _GEN_368; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_370 = 3'h1 == pht_rindex & 6'h32 == pht_raddr ? pht_1_50 : _GEN_369; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_371 = 3'h1 == pht_rindex & 6'h33 == pht_raddr ? pht_1_51 : _GEN_370; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_372 = 3'h1 == pht_rindex & 6'h34 == pht_raddr ? pht_1_52 : _GEN_371; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_373 = 3'h1 == pht_rindex & 6'h35 == pht_raddr ? pht_1_53 : _GEN_372; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_374 = 3'h1 == pht_rindex & 6'h36 == pht_raddr ? pht_1_54 : _GEN_373; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_375 = 3'h1 == pht_rindex & 6'h37 == pht_raddr ? pht_1_55 : _GEN_374; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_376 = 3'h1 == pht_rindex & 6'h38 == pht_raddr ? pht_1_56 : _GEN_375; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_377 = 3'h1 == pht_rindex & 6'h39 == pht_raddr ? pht_1_57 : _GEN_376; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_378 = 3'h1 == pht_rindex & 6'h3a == pht_raddr ? pht_1_58 : _GEN_377; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_379 = 3'h1 == pht_rindex & 6'h3b == pht_raddr ? pht_1_59 : _GEN_378; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_380 = 3'h1 == pht_rindex & 6'h3c == pht_raddr ? pht_1_60 : _GEN_379; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_381 = 3'h1 == pht_rindex & 6'h3d == pht_raddr ? pht_1_61 : _GEN_380; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_382 = 3'h1 == pht_rindex & 6'h3e == pht_raddr ? pht_1_62 : _GEN_381; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_383 = 3'h1 == pht_rindex & 6'h3f == pht_raddr ? pht_1_63 : _GEN_382; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_384 = 3'h1 == pht_rindex & 7'h40 == _GEN_9154 ? pht_1_64 : _GEN_383; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_385 = 3'h1 == pht_rindex & 7'h41 == _GEN_9154 ? pht_1_65 : _GEN_384; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_386 = 3'h1 == pht_rindex & 7'h42 == _GEN_9154 ? pht_1_66 : _GEN_385; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_387 = 3'h1 == pht_rindex & 7'h43 == _GEN_9154 ? pht_1_67 : _GEN_386; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_388 = 3'h1 == pht_rindex & 7'h44 == _GEN_9154 ? pht_1_68 : _GEN_387; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_389 = 3'h1 == pht_rindex & 7'h45 == _GEN_9154 ? pht_1_69 : _GEN_388; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_390 = 3'h1 == pht_rindex & 7'h46 == _GEN_9154 ? pht_1_70 : _GEN_389; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_391 = 3'h1 == pht_rindex & 7'h47 == _GEN_9154 ? pht_1_71 : _GEN_390; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_392 = 3'h1 == pht_rindex & 7'h48 == _GEN_9154 ? pht_1_72 : _GEN_391; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_393 = 3'h1 == pht_rindex & 7'h49 == _GEN_9154 ? pht_1_73 : _GEN_392; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_394 = 3'h1 == pht_rindex & 7'h4a == _GEN_9154 ? pht_1_74 : _GEN_393; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_395 = 3'h1 == pht_rindex & 7'h4b == _GEN_9154 ? pht_1_75 : _GEN_394; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_396 = 3'h1 == pht_rindex & 7'h4c == _GEN_9154 ? pht_1_76 : _GEN_395; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_397 = 3'h1 == pht_rindex & 7'h4d == _GEN_9154 ? pht_1_77 : _GEN_396; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_398 = 3'h1 == pht_rindex & 7'h4e == _GEN_9154 ? pht_1_78 : _GEN_397; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_399 = 3'h1 == pht_rindex & 7'h4f == _GEN_9154 ? pht_1_79 : _GEN_398; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_400 = 3'h1 == pht_rindex & 7'h50 == _GEN_9154 ? pht_1_80 : _GEN_399; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_401 = 3'h1 == pht_rindex & 7'h51 == _GEN_9154 ? pht_1_81 : _GEN_400; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_402 = 3'h1 == pht_rindex & 7'h52 == _GEN_9154 ? pht_1_82 : _GEN_401; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_403 = 3'h1 == pht_rindex & 7'h53 == _GEN_9154 ? pht_1_83 : _GEN_402; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_404 = 3'h1 == pht_rindex & 7'h54 == _GEN_9154 ? pht_1_84 : _GEN_403; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_405 = 3'h1 == pht_rindex & 7'h55 == _GEN_9154 ? pht_1_85 : _GEN_404; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_406 = 3'h1 == pht_rindex & 7'h56 == _GEN_9154 ? pht_1_86 : _GEN_405; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_407 = 3'h1 == pht_rindex & 7'h57 == _GEN_9154 ? pht_1_87 : _GEN_406; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_408 = 3'h1 == pht_rindex & 7'h58 == _GEN_9154 ? pht_1_88 : _GEN_407; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_409 = 3'h1 == pht_rindex & 7'h59 == _GEN_9154 ? pht_1_89 : _GEN_408; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_410 = 3'h1 == pht_rindex & 7'h5a == _GEN_9154 ? pht_1_90 : _GEN_409; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_411 = 3'h1 == pht_rindex & 7'h5b == _GEN_9154 ? pht_1_91 : _GEN_410; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_412 = 3'h1 == pht_rindex & 7'h5c == _GEN_9154 ? pht_1_92 : _GEN_411; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_413 = 3'h1 == pht_rindex & 7'h5d == _GEN_9154 ? pht_1_93 : _GEN_412; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_414 = 3'h1 == pht_rindex & 7'h5e == _GEN_9154 ? pht_1_94 : _GEN_413; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_415 = 3'h1 == pht_rindex & 7'h5f == _GEN_9154 ? pht_1_95 : _GEN_414; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_416 = 3'h1 == pht_rindex & 7'h60 == _GEN_9154 ? pht_1_96 : _GEN_415; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_417 = 3'h1 == pht_rindex & 7'h61 == _GEN_9154 ? pht_1_97 : _GEN_416; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_418 = 3'h1 == pht_rindex & 7'h62 == _GEN_9154 ? pht_1_98 : _GEN_417; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_419 = 3'h1 == pht_rindex & 7'h63 == _GEN_9154 ? pht_1_99 : _GEN_418; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_420 = 3'h1 == pht_rindex & 7'h64 == _GEN_9154 ? pht_1_100 : _GEN_419; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_421 = 3'h1 == pht_rindex & 7'h65 == _GEN_9154 ? pht_1_101 : _GEN_420; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_422 = 3'h1 == pht_rindex & 7'h66 == _GEN_9154 ? pht_1_102 : _GEN_421; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_423 = 3'h1 == pht_rindex & 7'h67 == _GEN_9154 ? pht_1_103 : _GEN_422; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_424 = 3'h1 == pht_rindex & 7'h68 == _GEN_9154 ? pht_1_104 : _GEN_423; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_425 = 3'h1 == pht_rindex & 7'h69 == _GEN_9154 ? pht_1_105 : _GEN_424; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_426 = 3'h1 == pht_rindex & 7'h6a == _GEN_9154 ? pht_1_106 : _GEN_425; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_427 = 3'h1 == pht_rindex & 7'h6b == _GEN_9154 ? pht_1_107 : _GEN_426; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_428 = 3'h1 == pht_rindex & 7'h6c == _GEN_9154 ? pht_1_108 : _GEN_427; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_429 = 3'h1 == pht_rindex & 7'h6d == _GEN_9154 ? pht_1_109 : _GEN_428; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_430 = 3'h1 == pht_rindex & 7'h6e == _GEN_9154 ? pht_1_110 : _GEN_429; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_431 = 3'h1 == pht_rindex & 7'h6f == _GEN_9154 ? pht_1_111 : _GEN_430; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_432 = 3'h1 == pht_rindex & 7'h70 == _GEN_9154 ? pht_1_112 : _GEN_431; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_433 = 3'h1 == pht_rindex & 7'h71 == _GEN_9154 ? pht_1_113 : _GEN_432; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_434 = 3'h1 == pht_rindex & 7'h72 == _GEN_9154 ? pht_1_114 : _GEN_433; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_435 = 3'h1 == pht_rindex & 7'h73 == _GEN_9154 ? pht_1_115 : _GEN_434; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_436 = 3'h1 == pht_rindex & 7'h74 == _GEN_9154 ? pht_1_116 : _GEN_435; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_437 = 3'h1 == pht_rindex & 7'h75 == _GEN_9154 ? pht_1_117 : _GEN_436; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_438 = 3'h1 == pht_rindex & 7'h76 == _GEN_9154 ? pht_1_118 : _GEN_437; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_439 = 3'h1 == pht_rindex & 7'h77 == _GEN_9154 ? pht_1_119 : _GEN_438; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_440 = 3'h1 == pht_rindex & 7'h78 == _GEN_9154 ? pht_1_120 : _GEN_439; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_441 = 3'h1 == pht_rindex & 7'h79 == _GEN_9154 ? pht_1_121 : _GEN_440; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_442 = 3'h1 == pht_rindex & 7'h7a == _GEN_9154 ? pht_1_122 : _GEN_441; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_443 = 3'h1 == pht_rindex & 7'h7b == _GEN_9154 ? pht_1_123 : _GEN_442; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_444 = 3'h1 == pht_rindex & 7'h7c == _GEN_9154 ? pht_1_124 : _GEN_443; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_445 = 3'h1 == pht_rindex & 7'h7d == _GEN_9154 ? pht_1_125 : _GEN_444; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_446 = 3'h1 == pht_rindex & 7'h7e == _GEN_9154 ? pht_1_126 : _GEN_445; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_447 = 3'h1 == pht_rindex & 7'h7f == _GEN_9154 ? pht_1_127 : _GEN_446; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_448 = 3'h1 == pht_rindex & 8'h80 == _GEN_9346 ? pht_1_128 : _GEN_447; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_449 = 3'h1 == pht_rindex & 8'h81 == _GEN_9346 ? pht_1_129 : _GEN_448; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_450 = 3'h1 == pht_rindex & 8'h82 == _GEN_9346 ? pht_1_130 : _GEN_449; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_451 = 3'h1 == pht_rindex & 8'h83 == _GEN_9346 ? pht_1_131 : _GEN_450; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_452 = 3'h1 == pht_rindex & 8'h84 == _GEN_9346 ? pht_1_132 : _GEN_451; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_453 = 3'h1 == pht_rindex & 8'h85 == _GEN_9346 ? pht_1_133 : _GEN_452; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_454 = 3'h1 == pht_rindex & 8'h86 == _GEN_9346 ? pht_1_134 : _GEN_453; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_455 = 3'h1 == pht_rindex & 8'h87 == _GEN_9346 ? pht_1_135 : _GEN_454; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_456 = 3'h1 == pht_rindex & 8'h88 == _GEN_9346 ? pht_1_136 : _GEN_455; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_457 = 3'h1 == pht_rindex & 8'h89 == _GEN_9346 ? pht_1_137 : _GEN_456; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_458 = 3'h1 == pht_rindex & 8'h8a == _GEN_9346 ? pht_1_138 : _GEN_457; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_459 = 3'h1 == pht_rindex & 8'h8b == _GEN_9346 ? pht_1_139 : _GEN_458; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_460 = 3'h1 == pht_rindex & 8'h8c == _GEN_9346 ? pht_1_140 : _GEN_459; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_461 = 3'h1 == pht_rindex & 8'h8d == _GEN_9346 ? pht_1_141 : _GEN_460; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_462 = 3'h1 == pht_rindex & 8'h8e == _GEN_9346 ? pht_1_142 : _GEN_461; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_463 = 3'h1 == pht_rindex & 8'h8f == _GEN_9346 ? pht_1_143 : _GEN_462; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_464 = 3'h1 == pht_rindex & 8'h90 == _GEN_9346 ? pht_1_144 : _GEN_463; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_465 = 3'h1 == pht_rindex & 8'h91 == _GEN_9346 ? pht_1_145 : _GEN_464; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_466 = 3'h1 == pht_rindex & 8'h92 == _GEN_9346 ? pht_1_146 : _GEN_465; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_467 = 3'h1 == pht_rindex & 8'h93 == _GEN_9346 ? pht_1_147 : _GEN_466; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_468 = 3'h1 == pht_rindex & 8'h94 == _GEN_9346 ? pht_1_148 : _GEN_467; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_469 = 3'h1 == pht_rindex & 8'h95 == _GEN_9346 ? pht_1_149 : _GEN_468; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_470 = 3'h1 == pht_rindex & 8'h96 == _GEN_9346 ? pht_1_150 : _GEN_469; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_471 = 3'h1 == pht_rindex & 8'h97 == _GEN_9346 ? pht_1_151 : _GEN_470; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_472 = 3'h1 == pht_rindex & 8'h98 == _GEN_9346 ? pht_1_152 : _GEN_471; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_473 = 3'h1 == pht_rindex & 8'h99 == _GEN_9346 ? pht_1_153 : _GEN_472; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_474 = 3'h1 == pht_rindex & 8'h9a == _GEN_9346 ? pht_1_154 : _GEN_473; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_475 = 3'h1 == pht_rindex & 8'h9b == _GEN_9346 ? pht_1_155 : _GEN_474; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_476 = 3'h1 == pht_rindex & 8'h9c == _GEN_9346 ? pht_1_156 : _GEN_475; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_477 = 3'h1 == pht_rindex & 8'h9d == _GEN_9346 ? pht_1_157 : _GEN_476; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_478 = 3'h1 == pht_rindex & 8'h9e == _GEN_9346 ? pht_1_158 : _GEN_477; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_479 = 3'h1 == pht_rindex & 8'h9f == _GEN_9346 ? pht_1_159 : _GEN_478; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_480 = 3'h1 == pht_rindex & 8'ha0 == _GEN_9346 ? pht_1_160 : _GEN_479; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_481 = 3'h1 == pht_rindex & 8'ha1 == _GEN_9346 ? pht_1_161 : _GEN_480; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_482 = 3'h1 == pht_rindex & 8'ha2 == _GEN_9346 ? pht_1_162 : _GEN_481; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_483 = 3'h1 == pht_rindex & 8'ha3 == _GEN_9346 ? pht_1_163 : _GEN_482; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_484 = 3'h1 == pht_rindex & 8'ha4 == _GEN_9346 ? pht_1_164 : _GEN_483; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_485 = 3'h1 == pht_rindex & 8'ha5 == _GEN_9346 ? pht_1_165 : _GEN_484; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_486 = 3'h1 == pht_rindex & 8'ha6 == _GEN_9346 ? pht_1_166 : _GEN_485; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_487 = 3'h1 == pht_rindex & 8'ha7 == _GEN_9346 ? pht_1_167 : _GEN_486; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_488 = 3'h1 == pht_rindex & 8'ha8 == _GEN_9346 ? pht_1_168 : _GEN_487; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_489 = 3'h1 == pht_rindex & 8'ha9 == _GEN_9346 ? pht_1_169 : _GEN_488; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_490 = 3'h1 == pht_rindex & 8'haa == _GEN_9346 ? pht_1_170 : _GEN_489; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_491 = 3'h1 == pht_rindex & 8'hab == _GEN_9346 ? pht_1_171 : _GEN_490; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_492 = 3'h1 == pht_rindex & 8'hac == _GEN_9346 ? pht_1_172 : _GEN_491; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_493 = 3'h1 == pht_rindex & 8'had == _GEN_9346 ? pht_1_173 : _GEN_492; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_494 = 3'h1 == pht_rindex & 8'hae == _GEN_9346 ? pht_1_174 : _GEN_493; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_495 = 3'h1 == pht_rindex & 8'haf == _GEN_9346 ? pht_1_175 : _GEN_494; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_496 = 3'h1 == pht_rindex & 8'hb0 == _GEN_9346 ? pht_1_176 : _GEN_495; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_497 = 3'h1 == pht_rindex & 8'hb1 == _GEN_9346 ? pht_1_177 : _GEN_496; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_498 = 3'h1 == pht_rindex & 8'hb2 == _GEN_9346 ? pht_1_178 : _GEN_497; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_499 = 3'h1 == pht_rindex & 8'hb3 == _GEN_9346 ? pht_1_179 : _GEN_498; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_500 = 3'h1 == pht_rindex & 8'hb4 == _GEN_9346 ? pht_1_180 : _GEN_499; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_501 = 3'h1 == pht_rindex & 8'hb5 == _GEN_9346 ? pht_1_181 : _GEN_500; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_502 = 3'h1 == pht_rindex & 8'hb6 == _GEN_9346 ? pht_1_182 : _GEN_501; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_503 = 3'h1 == pht_rindex & 8'hb7 == _GEN_9346 ? pht_1_183 : _GEN_502; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_504 = 3'h1 == pht_rindex & 8'hb8 == _GEN_9346 ? pht_1_184 : _GEN_503; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_505 = 3'h1 == pht_rindex & 8'hb9 == _GEN_9346 ? pht_1_185 : _GEN_504; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_506 = 3'h1 == pht_rindex & 8'hba == _GEN_9346 ? pht_1_186 : _GEN_505; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_507 = 3'h1 == pht_rindex & 8'hbb == _GEN_9346 ? pht_1_187 : _GEN_506; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_508 = 3'h1 == pht_rindex & 8'hbc == _GEN_9346 ? pht_1_188 : _GEN_507; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_509 = 3'h1 == pht_rindex & 8'hbd == _GEN_9346 ? pht_1_189 : _GEN_508; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_510 = 3'h1 == pht_rindex & 8'hbe == _GEN_9346 ? pht_1_190 : _GEN_509; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_511 = 3'h1 == pht_rindex & 8'hbf == _GEN_9346 ? pht_1_191 : _GEN_510; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_512 = 3'h1 == pht_rindex & 8'hc0 == _GEN_9346 ? pht_1_192 : _GEN_511; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_513 = 3'h1 == pht_rindex & 8'hc1 == _GEN_9346 ? pht_1_193 : _GEN_512; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_514 = 3'h1 == pht_rindex & 8'hc2 == _GEN_9346 ? pht_1_194 : _GEN_513; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_515 = 3'h1 == pht_rindex & 8'hc3 == _GEN_9346 ? pht_1_195 : _GEN_514; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_516 = 3'h1 == pht_rindex & 8'hc4 == _GEN_9346 ? pht_1_196 : _GEN_515; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_517 = 3'h1 == pht_rindex & 8'hc5 == _GEN_9346 ? pht_1_197 : _GEN_516; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_518 = 3'h1 == pht_rindex & 8'hc6 == _GEN_9346 ? pht_1_198 : _GEN_517; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_519 = 3'h1 == pht_rindex & 8'hc7 == _GEN_9346 ? pht_1_199 : _GEN_518; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_520 = 3'h1 == pht_rindex & 8'hc8 == _GEN_9346 ? pht_1_200 : _GEN_519; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_521 = 3'h1 == pht_rindex & 8'hc9 == _GEN_9346 ? pht_1_201 : _GEN_520; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_522 = 3'h1 == pht_rindex & 8'hca == _GEN_9346 ? pht_1_202 : _GEN_521; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_523 = 3'h1 == pht_rindex & 8'hcb == _GEN_9346 ? pht_1_203 : _GEN_522; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_524 = 3'h1 == pht_rindex & 8'hcc == _GEN_9346 ? pht_1_204 : _GEN_523; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_525 = 3'h1 == pht_rindex & 8'hcd == _GEN_9346 ? pht_1_205 : _GEN_524; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_526 = 3'h1 == pht_rindex & 8'hce == _GEN_9346 ? pht_1_206 : _GEN_525; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_527 = 3'h1 == pht_rindex & 8'hcf == _GEN_9346 ? pht_1_207 : _GEN_526; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_528 = 3'h1 == pht_rindex & 8'hd0 == _GEN_9346 ? pht_1_208 : _GEN_527; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_529 = 3'h1 == pht_rindex & 8'hd1 == _GEN_9346 ? pht_1_209 : _GEN_528; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_530 = 3'h1 == pht_rindex & 8'hd2 == _GEN_9346 ? pht_1_210 : _GEN_529; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_531 = 3'h1 == pht_rindex & 8'hd3 == _GEN_9346 ? pht_1_211 : _GEN_530; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_532 = 3'h1 == pht_rindex & 8'hd4 == _GEN_9346 ? pht_1_212 : _GEN_531; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_533 = 3'h1 == pht_rindex & 8'hd5 == _GEN_9346 ? pht_1_213 : _GEN_532; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_534 = 3'h1 == pht_rindex & 8'hd6 == _GEN_9346 ? pht_1_214 : _GEN_533; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_535 = 3'h1 == pht_rindex & 8'hd7 == _GEN_9346 ? pht_1_215 : _GEN_534; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_536 = 3'h1 == pht_rindex & 8'hd8 == _GEN_9346 ? pht_1_216 : _GEN_535; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_537 = 3'h1 == pht_rindex & 8'hd9 == _GEN_9346 ? pht_1_217 : _GEN_536; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_538 = 3'h1 == pht_rindex & 8'hda == _GEN_9346 ? pht_1_218 : _GEN_537; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_539 = 3'h1 == pht_rindex & 8'hdb == _GEN_9346 ? pht_1_219 : _GEN_538; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_540 = 3'h1 == pht_rindex & 8'hdc == _GEN_9346 ? pht_1_220 : _GEN_539; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_541 = 3'h1 == pht_rindex & 8'hdd == _GEN_9346 ? pht_1_221 : _GEN_540; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_542 = 3'h1 == pht_rindex & 8'hde == _GEN_9346 ? pht_1_222 : _GEN_541; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_543 = 3'h1 == pht_rindex & 8'hdf == _GEN_9346 ? pht_1_223 : _GEN_542; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_544 = 3'h1 == pht_rindex & 8'he0 == _GEN_9346 ? pht_1_224 : _GEN_543; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_545 = 3'h1 == pht_rindex & 8'he1 == _GEN_9346 ? pht_1_225 : _GEN_544; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_546 = 3'h1 == pht_rindex & 8'he2 == _GEN_9346 ? pht_1_226 : _GEN_545; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_547 = 3'h1 == pht_rindex & 8'he3 == _GEN_9346 ? pht_1_227 : _GEN_546; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_548 = 3'h1 == pht_rindex & 8'he4 == _GEN_9346 ? pht_1_228 : _GEN_547; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_549 = 3'h1 == pht_rindex & 8'he5 == _GEN_9346 ? pht_1_229 : _GEN_548; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_550 = 3'h1 == pht_rindex & 8'he6 == _GEN_9346 ? pht_1_230 : _GEN_549; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_551 = 3'h1 == pht_rindex & 8'he7 == _GEN_9346 ? pht_1_231 : _GEN_550; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_552 = 3'h1 == pht_rindex & 8'he8 == _GEN_9346 ? pht_1_232 : _GEN_551; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_553 = 3'h1 == pht_rindex & 8'he9 == _GEN_9346 ? pht_1_233 : _GEN_552; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_554 = 3'h1 == pht_rindex & 8'hea == _GEN_9346 ? pht_1_234 : _GEN_553; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_555 = 3'h1 == pht_rindex & 8'heb == _GEN_9346 ? pht_1_235 : _GEN_554; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_556 = 3'h1 == pht_rindex & 8'hec == _GEN_9346 ? pht_1_236 : _GEN_555; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_557 = 3'h1 == pht_rindex & 8'hed == _GEN_9346 ? pht_1_237 : _GEN_556; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_558 = 3'h1 == pht_rindex & 8'hee == _GEN_9346 ? pht_1_238 : _GEN_557; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_559 = 3'h1 == pht_rindex & 8'hef == _GEN_9346 ? pht_1_239 : _GEN_558; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_560 = 3'h1 == pht_rindex & 8'hf0 == _GEN_9346 ? pht_1_240 : _GEN_559; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_561 = 3'h1 == pht_rindex & 8'hf1 == _GEN_9346 ? pht_1_241 : _GEN_560; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_562 = 3'h1 == pht_rindex & 8'hf2 == _GEN_9346 ? pht_1_242 : _GEN_561; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_563 = 3'h1 == pht_rindex & 8'hf3 == _GEN_9346 ? pht_1_243 : _GEN_562; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_564 = 3'h1 == pht_rindex & 8'hf4 == _GEN_9346 ? pht_1_244 : _GEN_563; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_565 = 3'h1 == pht_rindex & 8'hf5 == _GEN_9346 ? pht_1_245 : _GEN_564; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_566 = 3'h1 == pht_rindex & 8'hf6 == _GEN_9346 ? pht_1_246 : _GEN_565; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_567 = 3'h1 == pht_rindex & 8'hf7 == _GEN_9346 ? pht_1_247 : _GEN_566; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_568 = 3'h1 == pht_rindex & 8'hf8 == _GEN_9346 ? pht_1_248 : _GEN_567; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_569 = 3'h1 == pht_rindex & 8'hf9 == _GEN_9346 ? pht_1_249 : _GEN_568; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_570 = 3'h1 == pht_rindex & 8'hfa == _GEN_9346 ? pht_1_250 : _GEN_569; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_571 = 3'h1 == pht_rindex & 8'hfb == _GEN_9346 ? pht_1_251 : _GEN_570; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_572 = 3'h1 == pht_rindex & 8'hfc == _GEN_9346 ? pht_1_252 : _GEN_571; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_573 = 3'h1 == pht_rindex & 8'hfd == _GEN_9346 ? pht_1_253 : _GEN_572; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_574 = 3'h1 == pht_rindex & 8'hfe == _GEN_9346 ? pht_1_254 : _GEN_573; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_575 = 3'h1 == pht_rindex & 8'hff == _GEN_9346 ? pht_1_255 : _GEN_574; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_576 = 3'h2 == pht_rindex & 6'h0 == pht_raddr ? pht_2_0 : _GEN_575; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_577 = 3'h2 == pht_rindex & 6'h1 == pht_raddr ? pht_2_1 : _GEN_576; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_578 = 3'h2 == pht_rindex & 6'h2 == pht_raddr ? pht_2_2 : _GEN_577; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_579 = 3'h2 == pht_rindex & 6'h3 == pht_raddr ? pht_2_3 : _GEN_578; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_580 = 3'h2 == pht_rindex & 6'h4 == pht_raddr ? pht_2_4 : _GEN_579; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_581 = 3'h2 == pht_rindex & 6'h5 == pht_raddr ? pht_2_5 : _GEN_580; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_582 = 3'h2 == pht_rindex & 6'h6 == pht_raddr ? pht_2_6 : _GEN_581; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_583 = 3'h2 == pht_rindex & 6'h7 == pht_raddr ? pht_2_7 : _GEN_582; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_584 = 3'h2 == pht_rindex & 6'h8 == pht_raddr ? pht_2_8 : _GEN_583; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_585 = 3'h2 == pht_rindex & 6'h9 == pht_raddr ? pht_2_9 : _GEN_584; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_586 = 3'h2 == pht_rindex & 6'ha == pht_raddr ? pht_2_10 : _GEN_585; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_587 = 3'h2 == pht_rindex & 6'hb == pht_raddr ? pht_2_11 : _GEN_586; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_588 = 3'h2 == pht_rindex & 6'hc == pht_raddr ? pht_2_12 : _GEN_587; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_589 = 3'h2 == pht_rindex & 6'hd == pht_raddr ? pht_2_13 : _GEN_588; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_590 = 3'h2 == pht_rindex & 6'he == pht_raddr ? pht_2_14 : _GEN_589; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_591 = 3'h2 == pht_rindex & 6'hf == pht_raddr ? pht_2_15 : _GEN_590; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_592 = 3'h2 == pht_rindex & 6'h10 == pht_raddr ? pht_2_16 : _GEN_591; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_593 = 3'h2 == pht_rindex & 6'h11 == pht_raddr ? pht_2_17 : _GEN_592; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_594 = 3'h2 == pht_rindex & 6'h12 == pht_raddr ? pht_2_18 : _GEN_593; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_595 = 3'h2 == pht_rindex & 6'h13 == pht_raddr ? pht_2_19 : _GEN_594; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_596 = 3'h2 == pht_rindex & 6'h14 == pht_raddr ? pht_2_20 : _GEN_595; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_597 = 3'h2 == pht_rindex & 6'h15 == pht_raddr ? pht_2_21 : _GEN_596; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_598 = 3'h2 == pht_rindex & 6'h16 == pht_raddr ? pht_2_22 : _GEN_597; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_599 = 3'h2 == pht_rindex & 6'h17 == pht_raddr ? pht_2_23 : _GEN_598; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_600 = 3'h2 == pht_rindex & 6'h18 == pht_raddr ? pht_2_24 : _GEN_599; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_601 = 3'h2 == pht_rindex & 6'h19 == pht_raddr ? pht_2_25 : _GEN_600; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_602 = 3'h2 == pht_rindex & 6'h1a == pht_raddr ? pht_2_26 : _GEN_601; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_603 = 3'h2 == pht_rindex & 6'h1b == pht_raddr ? pht_2_27 : _GEN_602; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_604 = 3'h2 == pht_rindex & 6'h1c == pht_raddr ? pht_2_28 : _GEN_603; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_605 = 3'h2 == pht_rindex & 6'h1d == pht_raddr ? pht_2_29 : _GEN_604; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_606 = 3'h2 == pht_rindex & 6'h1e == pht_raddr ? pht_2_30 : _GEN_605; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_607 = 3'h2 == pht_rindex & 6'h1f == pht_raddr ? pht_2_31 : _GEN_606; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_608 = 3'h2 == pht_rindex & 6'h20 == pht_raddr ? pht_2_32 : _GEN_607; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_609 = 3'h2 == pht_rindex & 6'h21 == pht_raddr ? pht_2_33 : _GEN_608; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_610 = 3'h2 == pht_rindex & 6'h22 == pht_raddr ? pht_2_34 : _GEN_609; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_611 = 3'h2 == pht_rindex & 6'h23 == pht_raddr ? pht_2_35 : _GEN_610; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_612 = 3'h2 == pht_rindex & 6'h24 == pht_raddr ? pht_2_36 : _GEN_611; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_613 = 3'h2 == pht_rindex & 6'h25 == pht_raddr ? pht_2_37 : _GEN_612; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_614 = 3'h2 == pht_rindex & 6'h26 == pht_raddr ? pht_2_38 : _GEN_613; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_615 = 3'h2 == pht_rindex & 6'h27 == pht_raddr ? pht_2_39 : _GEN_614; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_616 = 3'h2 == pht_rindex & 6'h28 == pht_raddr ? pht_2_40 : _GEN_615; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_617 = 3'h2 == pht_rindex & 6'h29 == pht_raddr ? pht_2_41 : _GEN_616; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_618 = 3'h2 == pht_rindex & 6'h2a == pht_raddr ? pht_2_42 : _GEN_617; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_619 = 3'h2 == pht_rindex & 6'h2b == pht_raddr ? pht_2_43 : _GEN_618; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_620 = 3'h2 == pht_rindex & 6'h2c == pht_raddr ? pht_2_44 : _GEN_619; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_621 = 3'h2 == pht_rindex & 6'h2d == pht_raddr ? pht_2_45 : _GEN_620; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_622 = 3'h2 == pht_rindex & 6'h2e == pht_raddr ? pht_2_46 : _GEN_621; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_623 = 3'h2 == pht_rindex & 6'h2f == pht_raddr ? pht_2_47 : _GEN_622; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_624 = 3'h2 == pht_rindex & 6'h30 == pht_raddr ? pht_2_48 : _GEN_623; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_625 = 3'h2 == pht_rindex & 6'h31 == pht_raddr ? pht_2_49 : _GEN_624; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_626 = 3'h2 == pht_rindex & 6'h32 == pht_raddr ? pht_2_50 : _GEN_625; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_627 = 3'h2 == pht_rindex & 6'h33 == pht_raddr ? pht_2_51 : _GEN_626; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_628 = 3'h2 == pht_rindex & 6'h34 == pht_raddr ? pht_2_52 : _GEN_627; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_629 = 3'h2 == pht_rindex & 6'h35 == pht_raddr ? pht_2_53 : _GEN_628; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_630 = 3'h2 == pht_rindex & 6'h36 == pht_raddr ? pht_2_54 : _GEN_629; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_631 = 3'h2 == pht_rindex & 6'h37 == pht_raddr ? pht_2_55 : _GEN_630; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_632 = 3'h2 == pht_rindex & 6'h38 == pht_raddr ? pht_2_56 : _GEN_631; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_633 = 3'h2 == pht_rindex & 6'h39 == pht_raddr ? pht_2_57 : _GEN_632; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_634 = 3'h2 == pht_rindex & 6'h3a == pht_raddr ? pht_2_58 : _GEN_633; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_635 = 3'h2 == pht_rindex & 6'h3b == pht_raddr ? pht_2_59 : _GEN_634; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_636 = 3'h2 == pht_rindex & 6'h3c == pht_raddr ? pht_2_60 : _GEN_635; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_637 = 3'h2 == pht_rindex & 6'h3d == pht_raddr ? pht_2_61 : _GEN_636; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_638 = 3'h2 == pht_rindex & 6'h3e == pht_raddr ? pht_2_62 : _GEN_637; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_639 = 3'h2 == pht_rindex & 6'h3f == pht_raddr ? pht_2_63 : _GEN_638; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_640 = 3'h2 == pht_rindex & 7'h40 == _GEN_9154 ? pht_2_64 : _GEN_639; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_641 = 3'h2 == pht_rindex & 7'h41 == _GEN_9154 ? pht_2_65 : _GEN_640; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_642 = 3'h2 == pht_rindex & 7'h42 == _GEN_9154 ? pht_2_66 : _GEN_641; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_643 = 3'h2 == pht_rindex & 7'h43 == _GEN_9154 ? pht_2_67 : _GEN_642; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_644 = 3'h2 == pht_rindex & 7'h44 == _GEN_9154 ? pht_2_68 : _GEN_643; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_645 = 3'h2 == pht_rindex & 7'h45 == _GEN_9154 ? pht_2_69 : _GEN_644; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_646 = 3'h2 == pht_rindex & 7'h46 == _GEN_9154 ? pht_2_70 : _GEN_645; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_647 = 3'h2 == pht_rindex & 7'h47 == _GEN_9154 ? pht_2_71 : _GEN_646; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_648 = 3'h2 == pht_rindex & 7'h48 == _GEN_9154 ? pht_2_72 : _GEN_647; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_649 = 3'h2 == pht_rindex & 7'h49 == _GEN_9154 ? pht_2_73 : _GEN_648; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_650 = 3'h2 == pht_rindex & 7'h4a == _GEN_9154 ? pht_2_74 : _GEN_649; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_651 = 3'h2 == pht_rindex & 7'h4b == _GEN_9154 ? pht_2_75 : _GEN_650; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_652 = 3'h2 == pht_rindex & 7'h4c == _GEN_9154 ? pht_2_76 : _GEN_651; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_653 = 3'h2 == pht_rindex & 7'h4d == _GEN_9154 ? pht_2_77 : _GEN_652; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_654 = 3'h2 == pht_rindex & 7'h4e == _GEN_9154 ? pht_2_78 : _GEN_653; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_655 = 3'h2 == pht_rindex & 7'h4f == _GEN_9154 ? pht_2_79 : _GEN_654; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_656 = 3'h2 == pht_rindex & 7'h50 == _GEN_9154 ? pht_2_80 : _GEN_655; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_657 = 3'h2 == pht_rindex & 7'h51 == _GEN_9154 ? pht_2_81 : _GEN_656; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_658 = 3'h2 == pht_rindex & 7'h52 == _GEN_9154 ? pht_2_82 : _GEN_657; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_659 = 3'h2 == pht_rindex & 7'h53 == _GEN_9154 ? pht_2_83 : _GEN_658; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_660 = 3'h2 == pht_rindex & 7'h54 == _GEN_9154 ? pht_2_84 : _GEN_659; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_661 = 3'h2 == pht_rindex & 7'h55 == _GEN_9154 ? pht_2_85 : _GEN_660; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_662 = 3'h2 == pht_rindex & 7'h56 == _GEN_9154 ? pht_2_86 : _GEN_661; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_663 = 3'h2 == pht_rindex & 7'h57 == _GEN_9154 ? pht_2_87 : _GEN_662; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_664 = 3'h2 == pht_rindex & 7'h58 == _GEN_9154 ? pht_2_88 : _GEN_663; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_665 = 3'h2 == pht_rindex & 7'h59 == _GEN_9154 ? pht_2_89 : _GEN_664; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_666 = 3'h2 == pht_rindex & 7'h5a == _GEN_9154 ? pht_2_90 : _GEN_665; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_667 = 3'h2 == pht_rindex & 7'h5b == _GEN_9154 ? pht_2_91 : _GEN_666; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_668 = 3'h2 == pht_rindex & 7'h5c == _GEN_9154 ? pht_2_92 : _GEN_667; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_669 = 3'h2 == pht_rindex & 7'h5d == _GEN_9154 ? pht_2_93 : _GEN_668; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_670 = 3'h2 == pht_rindex & 7'h5e == _GEN_9154 ? pht_2_94 : _GEN_669; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_671 = 3'h2 == pht_rindex & 7'h5f == _GEN_9154 ? pht_2_95 : _GEN_670; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_672 = 3'h2 == pht_rindex & 7'h60 == _GEN_9154 ? pht_2_96 : _GEN_671; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_673 = 3'h2 == pht_rindex & 7'h61 == _GEN_9154 ? pht_2_97 : _GEN_672; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_674 = 3'h2 == pht_rindex & 7'h62 == _GEN_9154 ? pht_2_98 : _GEN_673; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_675 = 3'h2 == pht_rindex & 7'h63 == _GEN_9154 ? pht_2_99 : _GEN_674; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_676 = 3'h2 == pht_rindex & 7'h64 == _GEN_9154 ? pht_2_100 : _GEN_675; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_677 = 3'h2 == pht_rindex & 7'h65 == _GEN_9154 ? pht_2_101 : _GEN_676; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_678 = 3'h2 == pht_rindex & 7'h66 == _GEN_9154 ? pht_2_102 : _GEN_677; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_679 = 3'h2 == pht_rindex & 7'h67 == _GEN_9154 ? pht_2_103 : _GEN_678; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_680 = 3'h2 == pht_rindex & 7'h68 == _GEN_9154 ? pht_2_104 : _GEN_679; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_681 = 3'h2 == pht_rindex & 7'h69 == _GEN_9154 ? pht_2_105 : _GEN_680; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_682 = 3'h2 == pht_rindex & 7'h6a == _GEN_9154 ? pht_2_106 : _GEN_681; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_683 = 3'h2 == pht_rindex & 7'h6b == _GEN_9154 ? pht_2_107 : _GEN_682; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_684 = 3'h2 == pht_rindex & 7'h6c == _GEN_9154 ? pht_2_108 : _GEN_683; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_685 = 3'h2 == pht_rindex & 7'h6d == _GEN_9154 ? pht_2_109 : _GEN_684; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_686 = 3'h2 == pht_rindex & 7'h6e == _GEN_9154 ? pht_2_110 : _GEN_685; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_687 = 3'h2 == pht_rindex & 7'h6f == _GEN_9154 ? pht_2_111 : _GEN_686; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_688 = 3'h2 == pht_rindex & 7'h70 == _GEN_9154 ? pht_2_112 : _GEN_687; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_689 = 3'h2 == pht_rindex & 7'h71 == _GEN_9154 ? pht_2_113 : _GEN_688; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_690 = 3'h2 == pht_rindex & 7'h72 == _GEN_9154 ? pht_2_114 : _GEN_689; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_691 = 3'h2 == pht_rindex & 7'h73 == _GEN_9154 ? pht_2_115 : _GEN_690; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_692 = 3'h2 == pht_rindex & 7'h74 == _GEN_9154 ? pht_2_116 : _GEN_691; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_693 = 3'h2 == pht_rindex & 7'h75 == _GEN_9154 ? pht_2_117 : _GEN_692; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_694 = 3'h2 == pht_rindex & 7'h76 == _GEN_9154 ? pht_2_118 : _GEN_693; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_695 = 3'h2 == pht_rindex & 7'h77 == _GEN_9154 ? pht_2_119 : _GEN_694; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_696 = 3'h2 == pht_rindex & 7'h78 == _GEN_9154 ? pht_2_120 : _GEN_695; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_697 = 3'h2 == pht_rindex & 7'h79 == _GEN_9154 ? pht_2_121 : _GEN_696; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_698 = 3'h2 == pht_rindex & 7'h7a == _GEN_9154 ? pht_2_122 : _GEN_697; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_699 = 3'h2 == pht_rindex & 7'h7b == _GEN_9154 ? pht_2_123 : _GEN_698; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_700 = 3'h2 == pht_rindex & 7'h7c == _GEN_9154 ? pht_2_124 : _GEN_699; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_701 = 3'h2 == pht_rindex & 7'h7d == _GEN_9154 ? pht_2_125 : _GEN_700; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_702 = 3'h2 == pht_rindex & 7'h7e == _GEN_9154 ? pht_2_126 : _GEN_701; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_703 = 3'h2 == pht_rindex & 7'h7f == _GEN_9154 ? pht_2_127 : _GEN_702; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_704 = 3'h2 == pht_rindex & 8'h80 == _GEN_9346 ? pht_2_128 : _GEN_703; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_705 = 3'h2 == pht_rindex & 8'h81 == _GEN_9346 ? pht_2_129 : _GEN_704; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_706 = 3'h2 == pht_rindex & 8'h82 == _GEN_9346 ? pht_2_130 : _GEN_705; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_707 = 3'h2 == pht_rindex & 8'h83 == _GEN_9346 ? pht_2_131 : _GEN_706; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_708 = 3'h2 == pht_rindex & 8'h84 == _GEN_9346 ? pht_2_132 : _GEN_707; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_709 = 3'h2 == pht_rindex & 8'h85 == _GEN_9346 ? pht_2_133 : _GEN_708; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_710 = 3'h2 == pht_rindex & 8'h86 == _GEN_9346 ? pht_2_134 : _GEN_709; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_711 = 3'h2 == pht_rindex & 8'h87 == _GEN_9346 ? pht_2_135 : _GEN_710; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_712 = 3'h2 == pht_rindex & 8'h88 == _GEN_9346 ? pht_2_136 : _GEN_711; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_713 = 3'h2 == pht_rindex & 8'h89 == _GEN_9346 ? pht_2_137 : _GEN_712; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_714 = 3'h2 == pht_rindex & 8'h8a == _GEN_9346 ? pht_2_138 : _GEN_713; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_715 = 3'h2 == pht_rindex & 8'h8b == _GEN_9346 ? pht_2_139 : _GEN_714; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_716 = 3'h2 == pht_rindex & 8'h8c == _GEN_9346 ? pht_2_140 : _GEN_715; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_717 = 3'h2 == pht_rindex & 8'h8d == _GEN_9346 ? pht_2_141 : _GEN_716; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_718 = 3'h2 == pht_rindex & 8'h8e == _GEN_9346 ? pht_2_142 : _GEN_717; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_719 = 3'h2 == pht_rindex & 8'h8f == _GEN_9346 ? pht_2_143 : _GEN_718; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_720 = 3'h2 == pht_rindex & 8'h90 == _GEN_9346 ? pht_2_144 : _GEN_719; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_721 = 3'h2 == pht_rindex & 8'h91 == _GEN_9346 ? pht_2_145 : _GEN_720; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_722 = 3'h2 == pht_rindex & 8'h92 == _GEN_9346 ? pht_2_146 : _GEN_721; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_723 = 3'h2 == pht_rindex & 8'h93 == _GEN_9346 ? pht_2_147 : _GEN_722; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_724 = 3'h2 == pht_rindex & 8'h94 == _GEN_9346 ? pht_2_148 : _GEN_723; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_725 = 3'h2 == pht_rindex & 8'h95 == _GEN_9346 ? pht_2_149 : _GEN_724; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_726 = 3'h2 == pht_rindex & 8'h96 == _GEN_9346 ? pht_2_150 : _GEN_725; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_727 = 3'h2 == pht_rindex & 8'h97 == _GEN_9346 ? pht_2_151 : _GEN_726; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_728 = 3'h2 == pht_rindex & 8'h98 == _GEN_9346 ? pht_2_152 : _GEN_727; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_729 = 3'h2 == pht_rindex & 8'h99 == _GEN_9346 ? pht_2_153 : _GEN_728; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_730 = 3'h2 == pht_rindex & 8'h9a == _GEN_9346 ? pht_2_154 : _GEN_729; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_731 = 3'h2 == pht_rindex & 8'h9b == _GEN_9346 ? pht_2_155 : _GEN_730; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_732 = 3'h2 == pht_rindex & 8'h9c == _GEN_9346 ? pht_2_156 : _GEN_731; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_733 = 3'h2 == pht_rindex & 8'h9d == _GEN_9346 ? pht_2_157 : _GEN_732; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_734 = 3'h2 == pht_rindex & 8'h9e == _GEN_9346 ? pht_2_158 : _GEN_733; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_735 = 3'h2 == pht_rindex & 8'h9f == _GEN_9346 ? pht_2_159 : _GEN_734; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_736 = 3'h2 == pht_rindex & 8'ha0 == _GEN_9346 ? pht_2_160 : _GEN_735; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_737 = 3'h2 == pht_rindex & 8'ha1 == _GEN_9346 ? pht_2_161 : _GEN_736; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_738 = 3'h2 == pht_rindex & 8'ha2 == _GEN_9346 ? pht_2_162 : _GEN_737; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_739 = 3'h2 == pht_rindex & 8'ha3 == _GEN_9346 ? pht_2_163 : _GEN_738; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_740 = 3'h2 == pht_rindex & 8'ha4 == _GEN_9346 ? pht_2_164 : _GEN_739; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_741 = 3'h2 == pht_rindex & 8'ha5 == _GEN_9346 ? pht_2_165 : _GEN_740; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_742 = 3'h2 == pht_rindex & 8'ha6 == _GEN_9346 ? pht_2_166 : _GEN_741; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_743 = 3'h2 == pht_rindex & 8'ha7 == _GEN_9346 ? pht_2_167 : _GEN_742; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_744 = 3'h2 == pht_rindex & 8'ha8 == _GEN_9346 ? pht_2_168 : _GEN_743; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_745 = 3'h2 == pht_rindex & 8'ha9 == _GEN_9346 ? pht_2_169 : _GEN_744; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_746 = 3'h2 == pht_rindex & 8'haa == _GEN_9346 ? pht_2_170 : _GEN_745; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_747 = 3'h2 == pht_rindex & 8'hab == _GEN_9346 ? pht_2_171 : _GEN_746; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_748 = 3'h2 == pht_rindex & 8'hac == _GEN_9346 ? pht_2_172 : _GEN_747; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_749 = 3'h2 == pht_rindex & 8'had == _GEN_9346 ? pht_2_173 : _GEN_748; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_750 = 3'h2 == pht_rindex & 8'hae == _GEN_9346 ? pht_2_174 : _GEN_749; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_751 = 3'h2 == pht_rindex & 8'haf == _GEN_9346 ? pht_2_175 : _GEN_750; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_752 = 3'h2 == pht_rindex & 8'hb0 == _GEN_9346 ? pht_2_176 : _GEN_751; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_753 = 3'h2 == pht_rindex & 8'hb1 == _GEN_9346 ? pht_2_177 : _GEN_752; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_754 = 3'h2 == pht_rindex & 8'hb2 == _GEN_9346 ? pht_2_178 : _GEN_753; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_755 = 3'h2 == pht_rindex & 8'hb3 == _GEN_9346 ? pht_2_179 : _GEN_754; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_756 = 3'h2 == pht_rindex & 8'hb4 == _GEN_9346 ? pht_2_180 : _GEN_755; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_757 = 3'h2 == pht_rindex & 8'hb5 == _GEN_9346 ? pht_2_181 : _GEN_756; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_758 = 3'h2 == pht_rindex & 8'hb6 == _GEN_9346 ? pht_2_182 : _GEN_757; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_759 = 3'h2 == pht_rindex & 8'hb7 == _GEN_9346 ? pht_2_183 : _GEN_758; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_760 = 3'h2 == pht_rindex & 8'hb8 == _GEN_9346 ? pht_2_184 : _GEN_759; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_761 = 3'h2 == pht_rindex & 8'hb9 == _GEN_9346 ? pht_2_185 : _GEN_760; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_762 = 3'h2 == pht_rindex & 8'hba == _GEN_9346 ? pht_2_186 : _GEN_761; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_763 = 3'h2 == pht_rindex & 8'hbb == _GEN_9346 ? pht_2_187 : _GEN_762; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_764 = 3'h2 == pht_rindex & 8'hbc == _GEN_9346 ? pht_2_188 : _GEN_763; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_765 = 3'h2 == pht_rindex & 8'hbd == _GEN_9346 ? pht_2_189 : _GEN_764; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_766 = 3'h2 == pht_rindex & 8'hbe == _GEN_9346 ? pht_2_190 : _GEN_765; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_767 = 3'h2 == pht_rindex & 8'hbf == _GEN_9346 ? pht_2_191 : _GEN_766; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_768 = 3'h2 == pht_rindex & 8'hc0 == _GEN_9346 ? pht_2_192 : _GEN_767; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_769 = 3'h2 == pht_rindex & 8'hc1 == _GEN_9346 ? pht_2_193 : _GEN_768; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_770 = 3'h2 == pht_rindex & 8'hc2 == _GEN_9346 ? pht_2_194 : _GEN_769; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_771 = 3'h2 == pht_rindex & 8'hc3 == _GEN_9346 ? pht_2_195 : _GEN_770; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_772 = 3'h2 == pht_rindex & 8'hc4 == _GEN_9346 ? pht_2_196 : _GEN_771; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_773 = 3'h2 == pht_rindex & 8'hc5 == _GEN_9346 ? pht_2_197 : _GEN_772; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_774 = 3'h2 == pht_rindex & 8'hc6 == _GEN_9346 ? pht_2_198 : _GEN_773; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_775 = 3'h2 == pht_rindex & 8'hc7 == _GEN_9346 ? pht_2_199 : _GEN_774; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_776 = 3'h2 == pht_rindex & 8'hc8 == _GEN_9346 ? pht_2_200 : _GEN_775; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_777 = 3'h2 == pht_rindex & 8'hc9 == _GEN_9346 ? pht_2_201 : _GEN_776; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_778 = 3'h2 == pht_rindex & 8'hca == _GEN_9346 ? pht_2_202 : _GEN_777; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_779 = 3'h2 == pht_rindex & 8'hcb == _GEN_9346 ? pht_2_203 : _GEN_778; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_780 = 3'h2 == pht_rindex & 8'hcc == _GEN_9346 ? pht_2_204 : _GEN_779; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_781 = 3'h2 == pht_rindex & 8'hcd == _GEN_9346 ? pht_2_205 : _GEN_780; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_782 = 3'h2 == pht_rindex & 8'hce == _GEN_9346 ? pht_2_206 : _GEN_781; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_783 = 3'h2 == pht_rindex & 8'hcf == _GEN_9346 ? pht_2_207 : _GEN_782; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_784 = 3'h2 == pht_rindex & 8'hd0 == _GEN_9346 ? pht_2_208 : _GEN_783; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_785 = 3'h2 == pht_rindex & 8'hd1 == _GEN_9346 ? pht_2_209 : _GEN_784; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_786 = 3'h2 == pht_rindex & 8'hd2 == _GEN_9346 ? pht_2_210 : _GEN_785; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_787 = 3'h2 == pht_rindex & 8'hd3 == _GEN_9346 ? pht_2_211 : _GEN_786; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_788 = 3'h2 == pht_rindex & 8'hd4 == _GEN_9346 ? pht_2_212 : _GEN_787; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_789 = 3'h2 == pht_rindex & 8'hd5 == _GEN_9346 ? pht_2_213 : _GEN_788; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_790 = 3'h2 == pht_rindex & 8'hd6 == _GEN_9346 ? pht_2_214 : _GEN_789; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_791 = 3'h2 == pht_rindex & 8'hd7 == _GEN_9346 ? pht_2_215 : _GEN_790; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_792 = 3'h2 == pht_rindex & 8'hd8 == _GEN_9346 ? pht_2_216 : _GEN_791; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_793 = 3'h2 == pht_rindex & 8'hd9 == _GEN_9346 ? pht_2_217 : _GEN_792; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_794 = 3'h2 == pht_rindex & 8'hda == _GEN_9346 ? pht_2_218 : _GEN_793; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_795 = 3'h2 == pht_rindex & 8'hdb == _GEN_9346 ? pht_2_219 : _GEN_794; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_796 = 3'h2 == pht_rindex & 8'hdc == _GEN_9346 ? pht_2_220 : _GEN_795; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_797 = 3'h2 == pht_rindex & 8'hdd == _GEN_9346 ? pht_2_221 : _GEN_796; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_798 = 3'h2 == pht_rindex & 8'hde == _GEN_9346 ? pht_2_222 : _GEN_797; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_799 = 3'h2 == pht_rindex & 8'hdf == _GEN_9346 ? pht_2_223 : _GEN_798; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_800 = 3'h2 == pht_rindex & 8'he0 == _GEN_9346 ? pht_2_224 : _GEN_799; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_801 = 3'h2 == pht_rindex & 8'he1 == _GEN_9346 ? pht_2_225 : _GEN_800; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_802 = 3'h2 == pht_rindex & 8'he2 == _GEN_9346 ? pht_2_226 : _GEN_801; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_803 = 3'h2 == pht_rindex & 8'he3 == _GEN_9346 ? pht_2_227 : _GEN_802; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_804 = 3'h2 == pht_rindex & 8'he4 == _GEN_9346 ? pht_2_228 : _GEN_803; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_805 = 3'h2 == pht_rindex & 8'he5 == _GEN_9346 ? pht_2_229 : _GEN_804; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_806 = 3'h2 == pht_rindex & 8'he6 == _GEN_9346 ? pht_2_230 : _GEN_805; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_807 = 3'h2 == pht_rindex & 8'he7 == _GEN_9346 ? pht_2_231 : _GEN_806; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_808 = 3'h2 == pht_rindex & 8'he8 == _GEN_9346 ? pht_2_232 : _GEN_807; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_809 = 3'h2 == pht_rindex & 8'he9 == _GEN_9346 ? pht_2_233 : _GEN_808; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_810 = 3'h2 == pht_rindex & 8'hea == _GEN_9346 ? pht_2_234 : _GEN_809; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_811 = 3'h2 == pht_rindex & 8'heb == _GEN_9346 ? pht_2_235 : _GEN_810; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_812 = 3'h2 == pht_rindex & 8'hec == _GEN_9346 ? pht_2_236 : _GEN_811; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_813 = 3'h2 == pht_rindex & 8'hed == _GEN_9346 ? pht_2_237 : _GEN_812; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_814 = 3'h2 == pht_rindex & 8'hee == _GEN_9346 ? pht_2_238 : _GEN_813; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_815 = 3'h2 == pht_rindex & 8'hef == _GEN_9346 ? pht_2_239 : _GEN_814; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_816 = 3'h2 == pht_rindex & 8'hf0 == _GEN_9346 ? pht_2_240 : _GEN_815; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_817 = 3'h2 == pht_rindex & 8'hf1 == _GEN_9346 ? pht_2_241 : _GEN_816; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_818 = 3'h2 == pht_rindex & 8'hf2 == _GEN_9346 ? pht_2_242 : _GEN_817; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_819 = 3'h2 == pht_rindex & 8'hf3 == _GEN_9346 ? pht_2_243 : _GEN_818; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_820 = 3'h2 == pht_rindex & 8'hf4 == _GEN_9346 ? pht_2_244 : _GEN_819; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_821 = 3'h2 == pht_rindex & 8'hf5 == _GEN_9346 ? pht_2_245 : _GEN_820; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_822 = 3'h2 == pht_rindex & 8'hf6 == _GEN_9346 ? pht_2_246 : _GEN_821; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_823 = 3'h2 == pht_rindex & 8'hf7 == _GEN_9346 ? pht_2_247 : _GEN_822; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_824 = 3'h2 == pht_rindex & 8'hf8 == _GEN_9346 ? pht_2_248 : _GEN_823; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_825 = 3'h2 == pht_rindex & 8'hf9 == _GEN_9346 ? pht_2_249 : _GEN_824; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_826 = 3'h2 == pht_rindex & 8'hfa == _GEN_9346 ? pht_2_250 : _GEN_825; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_827 = 3'h2 == pht_rindex & 8'hfb == _GEN_9346 ? pht_2_251 : _GEN_826; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_828 = 3'h2 == pht_rindex & 8'hfc == _GEN_9346 ? pht_2_252 : _GEN_827; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_829 = 3'h2 == pht_rindex & 8'hfd == _GEN_9346 ? pht_2_253 : _GEN_828; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_830 = 3'h2 == pht_rindex & 8'hfe == _GEN_9346 ? pht_2_254 : _GEN_829; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_831 = 3'h2 == pht_rindex & 8'hff == _GEN_9346 ? pht_2_255 : _GEN_830; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_832 = 3'h3 == pht_rindex & 6'h0 == pht_raddr ? pht_3_0 : _GEN_831; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_833 = 3'h3 == pht_rindex & 6'h1 == pht_raddr ? pht_3_1 : _GEN_832; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_834 = 3'h3 == pht_rindex & 6'h2 == pht_raddr ? pht_3_2 : _GEN_833; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_835 = 3'h3 == pht_rindex & 6'h3 == pht_raddr ? pht_3_3 : _GEN_834; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_836 = 3'h3 == pht_rindex & 6'h4 == pht_raddr ? pht_3_4 : _GEN_835; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_837 = 3'h3 == pht_rindex & 6'h5 == pht_raddr ? pht_3_5 : _GEN_836; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_838 = 3'h3 == pht_rindex & 6'h6 == pht_raddr ? pht_3_6 : _GEN_837; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_839 = 3'h3 == pht_rindex & 6'h7 == pht_raddr ? pht_3_7 : _GEN_838; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_840 = 3'h3 == pht_rindex & 6'h8 == pht_raddr ? pht_3_8 : _GEN_839; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_841 = 3'h3 == pht_rindex & 6'h9 == pht_raddr ? pht_3_9 : _GEN_840; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_842 = 3'h3 == pht_rindex & 6'ha == pht_raddr ? pht_3_10 : _GEN_841; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_843 = 3'h3 == pht_rindex & 6'hb == pht_raddr ? pht_3_11 : _GEN_842; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_844 = 3'h3 == pht_rindex & 6'hc == pht_raddr ? pht_3_12 : _GEN_843; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_845 = 3'h3 == pht_rindex & 6'hd == pht_raddr ? pht_3_13 : _GEN_844; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_846 = 3'h3 == pht_rindex & 6'he == pht_raddr ? pht_3_14 : _GEN_845; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_847 = 3'h3 == pht_rindex & 6'hf == pht_raddr ? pht_3_15 : _GEN_846; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_848 = 3'h3 == pht_rindex & 6'h10 == pht_raddr ? pht_3_16 : _GEN_847; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_849 = 3'h3 == pht_rindex & 6'h11 == pht_raddr ? pht_3_17 : _GEN_848; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_850 = 3'h3 == pht_rindex & 6'h12 == pht_raddr ? pht_3_18 : _GEN_849; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_851 = 3'h3 == pht_rindex & 6'h13 == pht_raddr ? pht_3_19 : _GEN_850; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_852 = 3'h3 == pht_rindex & 6'h14 == pht_raddr ? pht_3_20 : _GEN_851; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_853 = 3'h3 == pht_rindex & 6'h15 == pht_raddr ? pht_3_21 : _GEN_852; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_854 = 3'h3 == pht_rindex & 6'h16 == pht_raddr ? pht_3_22 : _GEN_853; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_855 = 3'h3 == pht_rindex & 6'h17 == pht_raddr ? pht_3_23 : _GEN_854; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_856 = 3'h3 == pht_rindex & 6'h18 == pht_raddr ? pht_3_24 : _GEN_855; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_857 = 3'h3 == pht_rindex & 6'h19 == pht_raddr ? pht_3_25 : _GEN_856; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_858 = 3'h3 == pht_rindex & 6'h1a == pht_raddr ? pht_3_26 : _GEN_857; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_859 = 3'h3 == pht_rindex & 6'h1b == pht_raddr ? pht_3_27 : _GEN_858; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_860 = 3'h3 == pht_rindex & 6'h1c == pht_raddr ? pht_3_28 : _GEN_859; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_861 = 3'h3 == pht_rindex & 6'h1d == pht_raddr ? pht_3_29 : _GEN_860; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_862 = 3'h3 == pht_rindex & 6'h1e == pht_raddr ? pht_3_30 : _GEN_861; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_863 = 3'h3 == pht_rindex & 6'h1f == pht_raddr ? pht_3_31 : _GEN_862; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_864 = 3'h3 == pht_rindex & 6'h20 == pht_raddr ? pht_3_32 : _GEN_863; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_865 = 3'h3 == pht_rindex & 6'h21 == pht_raddr ? pht_3_33 : _GEN_864; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_866 = 3'h3 == pht_rindex & 6'h22 == pht_raddr ? pht_3_34 : _GEN_865; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_867 = 3'h3 == pht_rindex & 6'h23 == pht_raddr ? pht_3_35 : _GEN_866; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_868 = 3'h3 == pht_rindex & 6'h24 == pht_raddr ? pht_3_36 : _GEN_867; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_869 = 3'h3 == pht_rindex & 6'h25 == pht_raddr ? pht_3_37 : _GEN_868; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_870 = 3'h3 == pht_rindex & 6'h26 == pht_raddr ? pht_3_38 : _GEN_869; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_871 = 3'h3 == pht_rindex & 6'h27 == pht_raddr ? pht_3_39 : _GEN_870; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_872 = 3'h3 == pht_rindex & 6'h28 == pht_raddr ? pht_3_40 : _GEN_871; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_873 = 3'h3 == pht_rindex & 6'h29 == pht_raddr ? pht_3_41 : _GEN_872; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_874 = 3'h3 == pht_rindex & 6'h2a == pht_raddr ? pht_3_42 : _GEN_873; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_875 = 3'h3 == pht_rindex & 6'h2b == pht_raddr ? pht_3_43 : _GEN_874; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_876 = 3'h3 == pht_rindex & 6'h2c == pht_raddr ? pht_3_44 : _GEN_875; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_877 = 3'h3 == pht_rindex & 6'h2d == pht_raddr ? pht_3_45 : _GEN_876; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_878 = 3'h3 == pht_rindex & 6'h2e == pht_raddr ? pht_3_46 : _GEN_877; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_879 = 3'h3 == pht_rindex & 6'h2f == pht_raddr ? pht_3_47 : _GEN_878; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_880 = 3'h3 == pht_rindex & 6'h30 == pht_raddr ? pht_3_48 : _GEN_879; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_881 = 3'h3 == pht_rindex & 6'h31 == pht_raddr ? pht_3_49 : _GEN_880; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_882 = 3'h3 == pht_rindex & 6'h32 == pht_raddr ? pht_3_50 : _GEN_881; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_883 = 3'h3 == pht_rindex & 6'h33 == pht_raddr ? pht_3_51 : _GEN_882; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_884 = 3'h3 == pht_rindex & 6'h34 == pht_raddr ? pht_3_52 : _GEN_883; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_885 = 3'h3 == pht_rindex & 6'h35 == pht_raddr ? pht_3_53 : _GEN_884; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_886 = 3'h3 == pht_rindex & 6'h36 == pht_raddr ? pht_3_54 : _GEN_885; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_887 = 3'h3 == pht_rindex & 6'h37 == pht_raddr ? pht_3_55 : _GEN_886; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_888 = 3'h3 == pht_rindex & 6'h38 == pht_raddr ? pht_3_56 : _GEN_887; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_889 = 3'h3 == pht_rindex & 6'h39 == pht_raddr ? pht_3_57 : _GEN_888; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_890 = 3'h3 == pht_rindex & 6'h3a == pht_raddr ? pht_3_58 : _GEN_889; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_891 = 3'h3 == pht_rindex & 6'h3b == pht_raddr ? pht_3_59 : _GEN_890; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_892 = 3'h3 == pht_rindex & 6'h3c == pht_raddr ? pht_3_60 : _GEN_891; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_893 = 3'h3 == pht_rindex & 6'h3d == pht_raddr ? pht_3_61 : _GEN_892; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_894 = 3'h3 == pht_rindex & 6'h3e == pht_raddr ? pht_3_62 : _GEN_893; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_895 = 3'h3 == pht_rindex & 6'h3f == pht_raddr ? pht_3_63 : _GEN_894; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_896 = 3'h3 == pht_rindex & 7'h40 == _GEN_9154 ? pht_3_64 : _GEN_895; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_897 = 3'h3 == pht_rindex & 7'h41 == _GEN_9154 ? pht_3_65 : _GEN_896; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_898 = 3'h3 == pht_rindex & 7'h42 == _GEN_9154 ? pht_3_66 : _GEN_897; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_899 = 3'h3 == pht_rindex & 7'h43 == _GEN_9154 ? pht_3_67 : _GEN_898; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_900 = 3'h3 == pht_rindex & 7'h44 == _GEN_9154 ? pht_3_68 : _GEN_899; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_901 = 3'h3 == pht_rindex & 7'h45 == _GEN_9154 ? pht_3_69 : _GEN_900; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_902 = 3'h3 == pht_rindex & 7'h46 == _GEN_9154 ? pht_3_70 : _GEN_901; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_903 = 3'h3 == pht_rindex & 7'h47 == _GEN_9154 ? pht_3_71 : _GEN_902; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_904 = 3'h3 == pht_rindex & 7'h48 == _GEN_9154 ? pht_3_72 : _GEN_903; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_905 = 3'h3 == pht_rindex & 7'h49 == _GEN_9154 ? pht_3_73 : _GEN_904; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_906 = 3'h3 == pht_rindex & 7'h4a == _GEN_9154 ? pht_3_74 : _GEN_905; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_907 = 3'h3 == pht_rindex & 7'h4b == _GEN_9154 ? pht_3_75 : _GEN_906; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_908 = 3'h3 == pht_rindex & 7'h4c == _GEN_9154 ? pht_3_76 : _GEN_907; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_909 = 3'h3 == pht_rindex & 7'h4d == _GEN_9154 ? pht_3_77 : _GEN_908; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_910 = 3'h3 == pht_rindex & 7'h4e == _GEN_9154 ? pht_3_78 : _GEN_909; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_911 = 3'h3 == pht_rindex & 7'h4f == _GEN_9154 ? pht_3_79 : _GEN_910; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_912 = 3'h3 == pht_rindex & 7'h50 == _GEN_9154 ? pht_3_80 : _GEN_911; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_913 = 3'h3 == pht_rindex & 7'h51 == _GEN_9154 ? pht_3_81 : _GEN_912; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_914 = 3'h3 == pht_rindex & 7'h52 == _GEN_9154 ? pht_3_82 : _GEN_913; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_915 = 3'h3 == pht_rindex & 7'h53 == _GEN_9154 ? pht_3_83 : _GEN_914; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_916 = 3'h3 == pht_rindex & 7'h54 == _GEN_9154 ? pht_3_84 : _GEN_915; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_917 = 3'h3 == pht_rindex & 7'h55 == _GEN_9154 ? pht_3_85 : _GEN_916; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_918 = 3'h3 == pht_rindex & 7'h56 == _GEN_9154 ? pht_3_86 : _GEN_917; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_919 = 3'h3 == pht_rindex & 7'h57 == _GEN_9154 ? pht_3_87 : _GEN_918; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_920 = 3'h3 == pht_rindex & 7'h58 == _GEN_9154 ? pht_3_88 : _GEN_919; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_921 = 3'h3 == pht_rindex & 7'h59 == _GEN_9154 ? pht_3_89 : _GEN_920; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_922 = 3'h3 == pht_rindex & 7'h5a == _GEN_9154 ? pht_3_90 : _GEN_921; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_923 = 3'h3 == pht_rindex & 7'h5b == _GEN_9154 ? pht_3_91 : _GEN_922; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_924 = 3'h3 == pht_rindex & 7'h5c == _GEN_9154 ? pht_3_92 : _GEN_923; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_925 = 3'h3 == pht_rindex & 7'h5d == _GEN_9154 ? pht_3_93 : _GEN_924; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_926 = 3'h3 == pht_rindex & 7'h5e == _GEN_9154 ? pht_3_94 : _GEN_925; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_927 = 3'h3 == pht_rindex & 7'h5f == _GEN_9154 ? pht_3_95 : _GEN_926; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_928 = 3'h3 == pht_rindex & 7'h60 == _GEN_9154 ? pht_3_96 : _GEN_927; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_929 = 3'h3 == pht_rindex & 7'h61 == _GEN_9154 ? pht_3_97 : _GEN_928; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_930 = 3'h3 == pht_rindex & 7'h62 == _GEN_9154 ? pht_3_98 : _GEN_929; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_931 = 3'h3 == pht_rindex & 7'h63 == _GEN_9154 ? pht_3_99 : _GEN_930; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_932 = 3'h3 == pht_rindex & 7'h64 == _GEN_9154 ? pht_3_100 : _GEN_931; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_933 = 3'h3 == pht_rindex & 7'h65 == _GEN_9154 ? pht_3_101 : _GEN_932; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_934 = 3'h3 == pht_rindex & 7'h66 == _GEN_9154 ? pht_3_102 : _GEN_933; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_935 = 3'h3 == pht_rindex & 7'h67 == _GEN_9154 ? pht_3_103 : _GEN_934; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_936 = 3'h3 == pht_rindex & 7'h68 == _GEN_9154 ? pht_3_104 : _GEN_935; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_937 = 3'h3 == pht_rindex & 7'h69 == _GEN_9154 ? pht_3_105 : _GEN_936; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_938 = 3'h3 == pht_rindex & 7'h6a == _GEN_9154 ? pht_3_106 : _GEN_937; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_939 = 3'h3 == pht_rindex & 7'h6b == _GEN_9154 ? pht_3_107 : _GEN_938; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_940 = 3'h3 == pht_rindex & 7'h6c == _GEN_9154 ? pht_3_108 : _GEN_939; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_941 = 3'h3 == pht_rindex & 7'h6d == _GEN_9154 ? pht_3_109 : _GEN_940; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_942 = 3'h3 == pht_rindex & 7'h6e == _GEN_9154 ? pht_3_110 : _GEN_941; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_943 = 3'h3 == pht_rindex & 7'h6f == _GEN_9154 ? pht_3_111 : _GEN_942; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_944 = 3'h3 == pht_rindex & 7'h70 == _GEN_9154 ? pht_3_112 : _GEN_943; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_945 = 3'h3 == pht_rindex & 7'h71 == _GEN_9154 ? pht_3_113 : _GEN_944; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_946 = 3'h3 == pht_rindex & 7'h72 == _GEN_9154 ? pht_3_114 : _GEN_945; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_947 = 3'h3 == pht_rindex & 7'h73 == _GEN_9154 ? pht_3_115 : _GEN_946; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_948 = 3'h3 == pht_rindex & 7'h74 == _GEN_9154 ? pht_3_116 : _GEN_947; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_949 = 3'h3 == pht_rindex & 7'h75 == _GEN_9154 ? pht_3_117 : _GEN_948; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_950 = 3'h3 == pht_rindex & 7'h76 == _GEN_9154 ? pht_3_118 : _GEN_949; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_951 = 3'h3 == pht_rindex & 7'h77 == _GEN_9154 ? pht_3_119 : _GEN_950; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_952 = 3'h3 == pht_rindex & 7'h78 == _GEN_9154 ? pht_3_120 : _GEN_951; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_953 = 3'h3 == pht_rindex & 7'h79 == _GEN_9154 ? pht_3_121 : _GEN_952; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_954 = 3'h3 == pht_rindex & 7'h7a == _GEN_9154 ? pht_3_122 : _GEN_953; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_955 = 3'h3 == pht_rindex & 7'h7b == _GEN_9154 ? pht_3_123 : _GEN_954; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_956 = 3'h3 == pht_rindex & 7'h7c == _GEN_9154 ? pht_3_124 : _GEN_955; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_957 = 3'h3 == pht_rindex & 7'h7d == _GEN_9154 ? pht_3_125 : _GEN_956; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_958 = 3'h3 == pht_rindex & 7'h7e == _GEN_9154 ? pht_3_126 : _GEN_957; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_959 = 3'h3 == pht_rindex & 7'h7f == _GEN_9154 ? pht_3_127 : _GEN_958; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_960 = 3'h3 == pht_rindex & 8'h80 == _GEN_9346 ? pht_3_128 : _GEN_959; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_961 = 3'h3 == pht_rindex & 8'h81 == _GEN_9346 ? pht_3_129 : _GEN_960; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_962 = 3'h3 == pht_rindex & 8'h82 == _GEN_9346 ? pht_3_130 : _GEN_961; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_963 = 3'h3 == pht_rindex & 8'h83 == _GEN_9346 ? pht_3_131 : _GEN_962; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_964 = 3'h3 == pht_rindex & 8'h84 == _GEN_9346 ? pht_3_132 : _GEN_963; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_965 = 3'h3 == pht_rindex & 8'h85 == _GEN_9346 ? pht_3_133 : _GEN_964; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_966 = 3'h3 == pht_rindex & 8'h86 == _GEN_9346 ? pht_3_134 : _GEN_965; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_967 = 3'h3 == pht_rindex & 8'h87 == _GEN_9346 ? pht_3_135 : _GEN_966; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_968 = 3'h3 == pht_rindex & 8'h88 == _GEN_9346 ? pht_3_136 : _GEN_967; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_969 = 3'h3 == pht_rindex & 8'h89 == _GEN_9346 ? pht_3_137 : _GEN_968; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_970 = 3'h3 == pht_rindex & 8'h8a == _GEN_9346 ? pht_3_138 : _GEN_969; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_971 = 3'h3 == pht_rindex & 8'h8b == _GEN_9346 ? pht_3_139 : _GEN_970; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_972 = 3'h3 == pht_rindex & 8'h8c == _GEN_9346 ? pht_3_140 : _GEN_971; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_973 = 3'h3 == pht_rindex & 8'h8d == _GEN_9346 ? pht_3_141 : _GEN_972; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_974 = 3'h3 == pht_rindex & 8'h8e == _GEN_9346 ? pht_3_142 : _GEN_973; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_975 = 3'h3 == pht_rindex & 8'h8f == _GEN_9346 ? pht_3_143 : _GEN_974; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_976 = 3'h3 == pht_rindex & 8'h90 == _GEN_9346 ? pht_3_144 : _GEN_975; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_977 = 3'h3 == pht_rindex & 8'h91 == _GEN_9346 ? pht_3_145 : _GEN_976; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_978 = 3'h3 == pht_rindex & 8'h92 == _GEN_9346 ? pht_3_146 : _GEN_977; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_979 = 3'h3 == pht_rindex & 8'h93 == _GEN_9346 ? pht_3_147 : _GEN_978; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_980 = 3'h3 == pht_rindex & 8'h94 == _GEN_9346 ? pht_3_148 : _GEN_979; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_981 = 3'h3 == pht_rindex & 8'h95 == _GEN_9346 ? pht_3_149 : _GEN_980; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_982 = 3'h3 == pht_rindex & 8'h96 == _GEN_9346 ? pht_3_150 : _GEN_981; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_983 = 3'h3 == pht_rindex & 8'h97 == _GEN_9346 ? pht_3_151 : _GEN_982; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_984 = 3'h3 == pht_rindex & 8'h98 == _GEN_9346 ? pht_3_152 : _GEN_983; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_985 = 3'h3 == pht_rindex & 8'h99 == _GEN_9346 ? pht_3_153 : _GEN_984; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_986 = 3'h3 == pht_rindex & 8'h9a == _GEN_9346 ? pht_3_154 : _GEN_985; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_987 = 3'h3 == pht_rindex & 8'h9b == _GEN_9346 ? pht_3_155 : _GEN_986; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_988 = 3'h3 == pht_rindex & 8'h9c == _GEN_9346 ? pht_3_156 : _GEN_987; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_989 = 3'h3 == pht_rindex & 8'h9d == _GEN_9346 ? pht_3_157 : _GEN_988; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_990 = 3'h3 == pht_rindex & 8'h9e == _GEN_9346 ? pht_3_158 : _GEN_989; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_991 = 3'h3 == pht_rindex & 8'h9f == _GEN_9346 ? pht_3_159 : _GEN_990; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_992 = 3'h3 == pht_rindex & 8'ha0 == _GEN_9346 ? pht_3_160 : _GEN_991; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_993 = 3'h3 == pht_rindex & 8'ha1 == _GEN_9346 ? pht_3_161 : _GEN_992; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_994 = 3'h3 == pht_rindex & 8'ha2 == _GEN_9346 ? pht_3_162 : _GEN_993; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_995 = 3'h3 == pht_rindex & 8'ha3 == _GEN_9346 ? pht_3_163 : _GEN_994; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_996 = 3'h3 == pht_rindex & 8'ha4 == _GEN_9346 ? pht_3_164 : _GEN_995; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_997 = 3'h3 == pht_rindex & 8'ha5 == _GEN_9346 ? pht_3_165 : _GEN_996; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_998 = 3'h3 == pht_rindex & 8'ha6 == _GEN_9346 ? pht_3_166 : _GEN_997; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_999 = 3'h3 == pht_rindex & 8'ha7 == _GEN_9346 ? pht_3_167 : _GEN_998; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1000 = 3'h3 == pht_rindex & 8'ha8 == _GEN_9346 ? pht_3_168 : _GEN_999; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1001 = 3'h3 == pht_rindex & 8'ha9 == _GEN_9346 ? pht_3_169 : _GEN_1000; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1002 = 3'h3 == pht_rindex & 8'haa == _GEN_9346 ? pht_3_170 : _GEN_1001; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1003 = 3'h3 == pht_rindex & 8'hab == _GEN_9346 ? pht_3_171 : _GEN_1002; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1004 = 3'h3 == pht_rindex & 8'hac == _GEN_9346 ? pht_3_172 : _GEN_1003; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1005 = 3'h3 == pht_rindex & 8'had == _GEN_9346 ? pht_3_173 : _GEN_1004; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1006 = 3'h3 == pht_rindex & 8'hae == _GEN_9346 ? pht_3_174 : _GEN_1005; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1007 = 3'h3 == pht_rindex & 8'haf == _GEN_9346 ? pht_3_175 : _GEN_1006; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1008 = 3'h3 == pht_rindex & 8'hb0 == _GEN_9346 ? pht_3_176 : _GEN_1007; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1009 = 3'h3 == pht_rindex & 8'hb1 == _GEN_9346 ? pht_3_177 : _GEN_1008; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1010 = 3'h3 == pht_rindex & 8'hb2 == _GEN_9346 ? pht_3_178 : _GEN_1009; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1011 = 3'h3 == pht_rindex & 8'hb3 == _GEN_9346 ? pht_3_179 : _GEN_1010; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1012 = 3'h3 == pht_rindex & 8'hb4 == _GEN_9346 ? pht_3_180 : _GEN_1011; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1013 = 3'h3 == pht_rindex & 8'hb5 == _GEN_9346 ? pht_3_181 : _GEN_1012; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1014 = 3'h3 == pht_rindex & 8'hb6 == _GEN_9346 ? pht_3_182 : _GEN_1013; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1015 = 3'h3 == pht_rindex & 8'hb7 == _GEN_9346 ? pht_3_183 : _GEN_1014; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1016 = 3'h3 == pht_rindex & 8'hb8 == _GEN_9346 ? pht_3_184 : _GEN_1015; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1017 = 3'h3 == pht_rindex & 8'hb9 == _GEN_9346 ? pht_3_185 : _GEN_1016; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1018 = 3'h3 == pht_rindex & 8'hba == _GEN_9346 ? pht_3_186 : _GEN_1017; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1019 = 3'h3 == pht_rindex & 8'hbb == _GEN_9346 ? pht_3_187 : _GEN_1018; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1020 = 3'h3 == pht_rindex & 8'hbc == _GEN_9346 ? pht_3_188 : _GEN_1019; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1021 = 3'h3 == pht_rindex & 8'hbd == _GEN_9346 ? pht_3_189 : _GEN_1020; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1022 = 3'h3 == pht_rindex & 8'hbe == _GEN_9346 ? pht_3_190 : _GEN_1021; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1023 = 3'h3 == pht_rindex & 8'hbf == _GEN_9346 ? pht_3_191 : _GEN_1022; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1024 = 3'h3 == pht_rindex & 8'hc0 == _GEN_9346 ? pht_3_192 : _GEN_1023; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1025 = 3'h3 == pht_rindex & 8'hc1 == _GEN_9346 ? pht_3_193 : _GEN_1024; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1026 = 3'h3 == pht_rindex & 8'hc2 == _GEN_9346 ? pht_3_194 : _GEN_1025; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1027 = 3'h3 == pht_rindex & 8'hc3 == _GEN_9346 ? pht_3_195 : _GEN_1026; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1028 = 3'h3 == pht_rindex & 8'hc4 == _GEN_9346 ? pht_3_196 : _GEN_1027; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1029 = 3'h3 == pht_rindex & 8'hc5 == _GEN_9346 ? pht_3_197 : _GEN_1028; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1030 = 3'h3 == pht_rindex & 8'hc6 == _GEN_9346 ? pht_3_198 : _GEN_1029; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1031 = 3'h3 == pht_rindex & 8'hc7 == _GEN_9346 ? pht_3_199 : _GEN_1030; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1032 = 3'h3 == pht_rindex & 8'hc8 == _GEN_9346 ? pht_3_200 : _GEN_1031; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1033 = 3'h3 == pht_rindex & 8'hc9 == _GEN_9346 ? pht_3_201 : _GEN_1032; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1034 = 3'h3 == pht_rindex & 8'hca == _GEN_9346 ? pht_3_202 : _GEN_1033; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1035 = 3'h3 == pht_rindex & 8'hcb == _GEN_9346 ? pht_3_203 : _GEN_1034; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1036 = 3'h3 == pht_rindex & 8'hcc == _GEN_9346 ? pht_3_204 : _GEN_1035; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1037 = 3'h3 == pht_rindex & 8'hcd == _GEN_9346 ? pht_3_205 : _GEN_1036; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1038 = 3'h3 == pht_rindex & 8'hce == _GEN_9346 ? pht_3_206 : _GEN_1037; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1039 = 3'h3 == pht_rindex & 8'hcf == _GEN_9346 ? pht_3_207 : _GEN_1038; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1040 = 3'h3 == pht_rindex & 8'hd0 == _GEN_9346 ? pht_3_208 : _GEN_1039; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1041 = 3'h3 == pht_rindex & 8'hd1 == _GEN_9346 ? pht_3_209 : _GEN_1040; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1042 = 3'h3 == pht_rindex & 8'hd2 == _GEN_9346 ? pht_3_210 : _GEN_1041; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1043 = 3'h3 == pht_rindex & 8'hd3 == _GEN_9346 ? pht_3_211 : _GEN_1042; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1044 = 3'h3 == pht_rindex & 8'hd4 == _GEN_9346 ? pht_3_212 : _GEN_1043; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1045 = 3'h3 == pht_rindex & 8'hd5 == _GEN_9346 ? pht_3_213 : _GEN_1044; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1046 = 3'h3 == pht_rindex & 8'hd6 == _GEN_9346 ? pht_3_214 : _GEN_1045; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1047 = 3'h3 == pht_rindex & 8'hd7 == _GEN_9346 ? pht_3_215 : _GEN_1046; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1048 = 3'h3 == pht_rindex & 8'hd8 == _GEN_9346 ? pht_3_216 : _GEN_1047; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1049 = 3'h3 == pht_rindex & 8'hd9 == _GEN_9346 ? pht_3_217 : _GEN_1048; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1050 = 3'h3 == pht_rindex & 8'hda == _GEN_9346 ? pht_3_218 : _GEN_1049; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1051 = 3'h3 == pht_rindex & 8'hdb == _GEN_9346 ? pht_3_219 : _GEN_1050; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1052 = 3'h3 == pht_rindex & 8'hdc == _GEN_9346 ? pht_3_220 : _GEN_1051; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1053 = 3'h3 == pht_rindex & 8'hdd == _GEN_9346 ? pht_3_221 : _GEN_1052; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1054 = 3'h3 == pht_rindex & 8'hde == _GEN_9346 ? pht_3_222 : _GEN_1053; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1055 = 3'h3 == pht_rindex & 8'hdf == _GEN_9346 ? pht_3_223 : _GEN_1054; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1056 = 3'h3 == pht_rindex & 8'he0 == _GEN_9346 ? pht_3_224 : _GEN_1055; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1057 = 3'h3 == pht_rindex & 8'he1 == _GEN_9346 ? pht_3_225 : _GEN_1056; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1058 = 3'h3 == pht_rindex & 8'he2 == _GEN_9346 ? pht_3_226 : _GEN_1057; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1059 = 3'h3 == pht_rindex & 8'he3 == _GEN_9346 ? pht_3_227 : _GEN_1058; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1060 = 3'h3 == pht_rindex & 8'he4 == _GEN_9346 ? pht_3_228 : _GEN_1059; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1061 = 3'h3 == pht_rindex & 8'he5 == _GEN_9346 ? pht_3_229 : _GEN_1060; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1062 = 3'h3 == pht_rindex & 8'he6 == _GEN_9346 ? pht_3_230 : _GEN_1061; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1063 = 3'h3 == pht_rindex & 8'he7 == _GEN_9346 ? pht_3_231 : _GEN_1062; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1064 = 3'h3 == pht_rindex & 8'he8 == _GEN_9346 ? pht_3_232 : _GEN_1063; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1065 = 3'h3 == pht_rindex & 8'he9 == _GEN_9346 ? pht_3_233 : _GEN_1064; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1066 = 3'h3 == pht_rindex & 8'hea == _GEN_9346 ? pht_3_234 : _GEN_1065; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1067 = 3'h3 == pht_rindex & 8'heb == _GEN_9346 ? pht_3_235 : _GEN_1066; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1068 = 3'h3 == pht_rindex & 8'hec == _GEN_9346 ? pht_3_236 : _GEN_1067; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1069 = 3'h3 == pht_rindex & 8'hed == _GEN_9346 ? pht_3_237 : _GEN_1068; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1070 = 3'h3 == pht_rindex & 8'hee == _GEN_9346 ? pht_3_238 : _GEN_1069; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1071 = 3'h3 == pht_rindex & 8'hef == _GEN_9346 ? pht_3_239 : _GEN_1070; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1072 = 3'h3 == pht_rindex & 8'hf0 == _GEN_9346 ? pht_3_240 : _GEN_1071; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1073 = 3'h3 == pht_rindex & 8'hf1 == _GEN_9346 ? pht_3_241 : _GEN_1072; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1074 = 3'h3 == pht_rindex & 8'hf2 == _GEN_9346 ? pht_3_242 : _GEN_1073; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1075 = 3'h3 == pht_rindex & 8'hf3 == _GEN_9346 ? pht_3_243 : _GEN_1074; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1076 = 3'h3 == pht_rindex & 8'hf4 == _GEN_9346 ? pht_3_244 : _GEN_1075; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1077 = 3'h3 == pht_rindex & 8'hf5 == _GEN_9346 ? pht_3_245 : _GEN_1076; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1078 = 3'h3 == pht_rindex & 8'hf6 == _GEN_9346 ? pht_3_246 : _GEN_1077; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1079 = 3'h3 == pht_rindex & 8'hf7 == _GEN_9346 ? pht_3_247 : _GEN_1078; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1080 = 3'h3 == pht_rindex & 8'hf8 == _GEN_9346 ? pht_3_248 : _GEN_1079; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1081 = 3'h3 == pht_rindex & 8'hf9 == _GEN_9346 ? pht_3_249 : _GEN_1080; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1082 = 3'h3 == pht_rindex & 8'hfa == _GEN_9346 ? pht_3_250 : _GEN_1081; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1083 = 3'h3 == pht_rindex & 8'hfb == _GEN_9346 ? pht_3_251 : _GEN_1082; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1084 = 3'h3 == pht_rindex & 8'hfc == _GEN_9346 ? pht_3_252 : _GEN_1083; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1085 = 3'h3 == pht_rindex & 8'hfd == _GEN_9346 ? pht_3_253 : _GEN_1084; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1086 = 3'h3 == pht_rindex & 8'hfe == _GEN_9346 ? pht_3_254 : _GEN_1085; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1087 = 3'h3 == pht_rindex & 8'hff == _GEN_9346 ? pht_3_255 : _GEN_1086; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1088 = 3'h4 == pht_rindex & 6'h0 == pht_raddr ? pht_4_0 : _GEN_1087; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1089 = 3'h4 == pht_rindex & 6'h1 == pht_raddr ? pht_4_1 : _GEN_1088; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1090 = 3'h4 == pht_rindex & 6'h2 == pht_raddr ? pht_4_2 : _GEN_1089; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1091 = 3'h4 == pht_rindex & 6'h3 == pht_raddr ? pht_4_3 : _GEN_1090; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1092 = 3'h4 == pht_rindex & 6'h4 == pht_raddr ? pht_4_4 : _GEN_1091; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1093 = 3'h4 == pht_rindex & 6'h5 == pht_raddr ? pht_4_5 : _GEN_1092; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1094 = 3'h4 == pht_rindex & 6'h6 == pht_raddr ? pht_4_6 : _GEN_1093; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1095 = 3'h4 == pht_rindex & 6'h7 == pht_raddr ? pht_4_7 : _GEN_1094; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1096 = 3'h4 == pht_rindex & 6'h8 == pht_raddr ? pht_4_8 : _GEN_1095; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1097 = 3'h4 == pht_rindex & 6'h9 == pht_raddr ? pht_4_9 : _GEN_1096; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1098 = 3'h4 == pht_rindex & 6'ha == pht_raddr ? pht_4_10 : _GEN_1097; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1099 = 3'h4 == pht_rindex & 6'hb == pht_raddr ? pht_4_11 : _GEN_1098; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1100 = 3'h4 == pht_rindex & 6'hc == pht_raddr ? pht_4_12 : _GEN_1099; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1101 = 3'h4 == pht_rindex & 6'hd == pht_raddr ? pht_4_13 : _GEN_1100; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1102 = 3'h4 == pht_rindex & 6'he == pht_raddr ? pht_4_14 : _GEN_1101; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1103 = 3'h4 == pht_rindex & 6'hf == pht_raddr ? pht_4_15 : _GEN_1102; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1104 = 3'h4 == pht_rindex & 6'h10 == pht_raddr ? pht_4_16 : _GEN_1103; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1105 = 3'h4 == pht_rindex & 6'h11 == pht_raddr ? pht_4_17 : _GEN_1104; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1106 = 3'h4 == pht_rindex & 6'h12 == pht_raddr ? pht_4_18 : _GEN_1105; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1107 = 3'h4 == pht_rindex & 6'h13 == pht_raddr ? pht_4_19 : _GEN_1106; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1108 = 3'h4 == pht_rindex & 6'h14 == pht_raddr ? pht_4_20 : _GEN_1107; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1109 = 3'h4 == pht_rindex & 6'h15 == pht_raddr ? pht_4_21 : _GEN_1108; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1110 = 3'h4 == pht_rindex & 6'h16 == pht_raddr ? pht_4_22 : _GEN_1109; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1111 = 3'h4 == pht_rindex & 6'h17 == pht_raddr ? pht_4_23 : _GEN_1110; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1112 = 3'h4 == pht_rindex & 6'h18 == pht_raddr ? pht_4_24 : _GEN_1111; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1113 = 3'h4 == pht_rindex & 6'h19 == pht_raddr ? pht_4_25 : _GEN_1112; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1114 = 3'h4 == pht_rindex & 6'h1a == pht_raddr ? pht_4_26 : _GEN_1113; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1115 = 3'h4 == pht_rindex & 6'h1b == pht_raddr ? pht_4_27 : _GEN_1114; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1116 = 3'h4 == pht_rindex & 6'h1c == pht_raddr ? pht_4_28 : _GEN_1115; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1117 = 3'h4 == pht_rindex & 6'h1d == pht_raddr ? pht_4_29 : _GEN_1116; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1118 = 3'h4 == pht_rindex & 6'h1e == pht_raddr ? pht_4_30 : _GEN_1117; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1119 = 3'h4 == pht_rindex & 6'h1f == pht_raddr ? pht_4_31 : _GEN_1118; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1120 = 3'h4 == pht_rindex & 6'h20 == pht_raddr ? pht_4_32 : _GEN_1119; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1121 = 3'h4 == pht_rindex & 6'h21 == pht_raddr ? pht_4_33 : _GEN_1120; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1122 = 3'h4 == pht_rindex & 6'h22 == pht_raddr ? pht_4_34 : _GEN_1121; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1123 = 3'h4 == pht_rindex & 6'h23 == pht_raddr ? pht_4_35 : _GEN_1122; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1124 = 3'h4 == pht_rindex & 6'h24 == pht_raddr ? pht_4_36 : _GEN_1123; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1125 = 3'h4 == pht_rindex & 6'h25 == pht_raddr ? pht_4_37 : _GEN_1124; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1126 = 3'h4 == pht_rindex & 6'h26 == pht_raddr ? pht_4_38 : _GEN_1125; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1127 = 3'h4 == pht_rindex & 6'h27 == pht_raddr ? pht_4_39 : _GEN_1126; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1128 = 3'h4 == pht_rindex & 6'h28 == pht_raddr ? pht_4_40 : _GEN_1127; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1129 = 3'h4 == pht_rindex & 6'h29 == pht_raddr ? pht_4_41 : _GEN_1128; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1130 = 3'h4 == pht_rindex & 6'h2a == pht_raddr ? pht_4_42 : _GEN_1129; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1131 = 3'h4 == pht_rindex & 6'h2b == pht_raddr ? pht_4_43 : _GEN_1130; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1132 = 3'h4 == pht_rindex & 6'h2c == pht_raddr ? pht_4_44 : _GEN_1131; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1133 = 3'h4 == pht_rindex & 6'h2d == pht_raddr ? pht_4_45 : _GEN_1132; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1134 = 3'h4 == pht_rindex & 6'h2e == pht_raddr ? pht_4_46 : _GEN_1133; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1135 = 3'h4 == pht_rindex & 6'h2f == pht_raddr ? pht_4_47 : _GEN_1134; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1136 = 3'h4 == pht_rindex & 6'h30 == pht_raddr ? pht_4_48 : _GEN_1135; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1137 = 3'h4 == pht_rindex & 6'h31 == pht_raddr ? pht_4_49 : _GEN_1136; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1138 = 3'h4 == pht_rindex & 6'h32 == pht_raddr ? pht_4_50 : _GEN_1137; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1139 = 3'h4 == pht_rindex & 6'h33 == pht_raddr ? pht_4_51 : _GEN_1138; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1140 = 3'h4 == pht_rindex & 6'h34 == pht_raddr ? pht_4_52 : _GEN_1139; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1141 = 3'h4 == pht_rindex & 6'h35 == pht_raddr ? pht_4_53 : _GEN_1140; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1142 = 3'h4 == pht_rindex & 6'h36 == pht_raddr ? pht_4_54 : _GEN_1141; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1143 = 3'h4 == pht_rindex & 6'h37 == pht_raddr ? pht_4_55 : _GEN_1142; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1144 = 3'h4 == pht_rindex & 6'h38 == pht_raddr ? pht_4_56 : _GEN_1143; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1145 = 3'h4 == pht_rindex & 6'h39 == pht_raddr ? pht_4_57 : _GEN_1144; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1146 = 3'h4 == pht_rindex & 6'h3a == pht_raddr ? pht_4_58 : _GEN_1145; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1147 = 3'h4 == pht_rindex & 6'h3b == pht_raddr ? pht_4_59 : _GEN_1146; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1148 = 3'h4 == pht_rindex & 6'h3c == pht_raddr ? pht_4_60 : _GEN_1147; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1149 = 3'h4 == pht_rindex & 6'h3d == pht_raddr ? pht_4_61 : _GEN_1148; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1150 = 3'h4 == pht_rindex & 6'h3e == pht_raddr ? pht_4_62 : _GEN_1149; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1151 = 3'h4 == pht_rindex & 6'h3f == pht_raddr ? pht_4_63 : _GEN_1150; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1152 = 3'h4 == pht_rindex & 7'h40 == _GEN_9154 ? pht_4_64 : _GEN_1151; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1153 = 3'h4 == pht_rindex & 7'h41 == _GEN_9154 ? pht_4_65 : _GEN_1152; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1154 = 3'h4 == pht_rindex & 7'h42 == _GEN_9154 ? pht_4_66 : _GEN_1153; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1155 = 3'h4 == pht_rindex & 7'h43 == _GEN_9154 ? pht_4_67 : _GEN_1154; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1156 = 3'h4 == pht_rindex & 7'h44 == _GEN_9154 ? pht_4_68 : _GEN_1155; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1157 = 3'h4 == pht_rindex & 7'h45 == _GEN_9154 ? pht_4_69 : _GEN_1156; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1158 = 3'h4 == pht_rindex & 7'h46 == _GEN_9154 ? pht_4_70 : _GEN_1157; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1159 = 3'h4 == pht_rindex & 7'h47 == _GEN_9154 ? pht_4_71 : _GEN_1158; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1160 = 3'h4 == pht_rindex & 7'h48 == _GEN_9154 ? pht_4_72 : _GEN_1159; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1161 = 3'h4 == pht_rindex & 7'h49 == _GEN_9154 ? pht_4_73 : _GEN_1160; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1162 = 3'h4 == pht_rindex & 7'h4a == _GEN_9154 ? pht_4_74 : _GEN_1161; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1163 = 3'h4 == pht_rindex & 7'h4b == _GEN_9154 ? pht_4_75 : _GEN_1162; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1164 = 3'h4 == pht_rindex & 7'h4c == _GEN_9154 ? pht_4_76 : _GEN_1163; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1165 = 3'h4 == pht_rindex & 7'h4d == _GEN_9154 ? pht_4_77 : _GEN_1164; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1166 = 3'h4 == pht_rindex & 7'h4e == _GEN_9154 ? pht_4_78 : _GEN_1165; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1167 = 3'h4 == pht_rindex & 7'h4f == _GEN_9154 ? pht_4_79 : _GEN_1166; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1168 = 3'h4 == pht_rindex & 7'h50 == _GEN_9154 ? pht_4_80 : _GEN_1167; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1169 = 3'h4 == pht_rindex & 7'h51 == _GEN_9154 ? pht_4_81 : _GEN_1168; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1170 = 3'h4 == pht_rindex & 7'h52 == _GEN_9154 ? pht_4_82 : _GEN_1169; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1171 = 3'h4 == pht_rindex & 7'h53 == _GEN_9154 ? pht_4_83 : _GEN_1170; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1172 = 3'h4 == pht_rindex & 7'h54 == _GEN_9154 ? pht_4_84 : _GEN_1171; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1173 = 3'h4 == pht_rindex & 7'h55 == _GEN_9154 ? pht_4_85 : _GEN_1172; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1174 = 3'h4 == pht_rindex & 7'h56 == _GEN_9154 ? pht_4_86 : _GEN_1173; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1175 = 3'h4 == pht_rindex & 7'h57 == _GEN_9154 ? pht_4_87 : _GEN_1174; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1176 = 3'h4 == pht_rindex & 7'h58 == _GEN_9154 ? pht_4_88 : _GEN_1175; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1177 = 3'h4 == pht_rindex & 7'h59 == _GEN_9154 ? pht_4_89 : _GEN_1176; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1178 = 3'h4 == pht_rindex & 7'h5a == _GEN_9154 ? pht_4_90 : _GEN_1177; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1179 = 3'h4 == pht_rindex & 7'h5b == _GEN_9154 ? pht_4_91 : _GEN_1178; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1180 = 3'h4 == pht_rindex & 7'h5c == _GEN_9154 ? pht_4_92 : _GEN_1179; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1181 = 3'h4 == pht_rindex & 7'h5d == _GEN_9154 ? pht_4_93 : _GEN_1180; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1182 = 3'h4 == pht_rindex & 7'h5e == _GEN_9154 ? pht_4_94 : _GEN_1181; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1183 = 3'h4 == pht_rindex & 7'h5f == _GEN_9154 ? pht_4_95 : _GEN_1182; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1184 = 3'h4 == pht_rindex & 7'h60 == _GEN_9154 ? pht_4_96 : _GEN_1183; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1185 = 3'h4 == pht_rindex & 7'h61 == _GEN_9154 ? pht_4_97 : _GEN_1184; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1186 = 3'h4 == pht_rindex & 7'h62 == _GEN_9154 ? pht_4_98 : _GEN_1185; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1187 = 3'h4 == pht_rindex & 7'h63 == _GEN_9154 ? pht_4_99 : _GEN_1186; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1188 = 3'h4 == pht_rindex & 7'h64 == _GEN_9154 ? pht_4_100 : _GEN_1187; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1189 = 3'h4 == pht_rindex & 7'h65 == _GEN_9154 ? pht_4_101 : _GEN_1188; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1190 = 3'h4 == pht_rindex & 7'h66 == _GEN_9154 ? pht_4_102 : _GEN_1189; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1191 = 3'h4 == pht_rindex & 7'h67 == _GEN_9154 ? pht_4_103 : _GEN_1190; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1192 = 3'h4 == pht_rindex & 7'h68 == _GEN_9154 ? pht_4_104 : _GEN_1191; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1193 = 3'h4 == pht_rindex & 7'h69 == _GEN_9154 ? pht_4_105 : _GEN_1192; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1194 = 3'h4 == pht_rindex & 7'h6a == _GEN_9154 ? pht_4_106 : _GEN_1193; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1195 = 3'h4 == pht_rindex & 7'h6b == _GEN_9154 ? pht_4_107 : _GEN_1194; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1196 = 3'h4 == pht_rindex & 7'h6c == _GEN_9154 ? pht_4_108 : _GEN_1195; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1197 = 3'h4 == pht_rindex & 7'h6d == _GEN_9154 ? pht_4_109 : _GEN_1196; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1198 = 3'h4 == pht_rindex & 7'h6e == _GEN_9154 ? pht_4_110 : _GEN_1197; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1199 = 3'h4 == pht_rindex & 7'h6f == _GEN_9154 ? pht_4_111 : _GEN_1198; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1200 = 3'h4 == pht_rindex & 7'h70 == _GEN_9154 ? pht_4_112 : _GEN_1199; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1201 = 3'h4 == pht_rindex & 7'h71 == _GEN_9154 ? pht_4_113 : _GEN_1200; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1202 = 3'h4 == pht_rindex & 7'h72 == _GEN_9154 ? pht_4_114 : _GEN_1201; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1203 = 3'h4 == pht_rindex & 7'h73 == _GEN_9154 ? pht_4_115 : _GEN_1202; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1204 = 3'h4 == pht_rindex & 7'h74 == _GEN_9154 ? pht_4_116 : _GEN_1203; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1205 = 3'h4 == pht_rindex & 7'h75 == _GEN_9154 ? pht_4_117 : _GEN_1204; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1206 = 3'h4 == pht_rindex & 7'h76 == _GEN_9154 ? pht_4_118 : _GEN_1205; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1207 = 3'h4 == pht_rindex & 7'h77 == _GEN_9154 ? pht_4_119 : _GEN_1206; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1208 = 3'h4 == pht_rindex & 7'h78 == _GEN_9154 ? pht_4_120 : _GEN_1207; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1209 = 3'h4 == pht_rindex & 7'h79 == _GEN_9154 ? pht_4_121 : _GEN_1208; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1210 = 3'h4 == pht_rindex & 7'h7a == _GEN_9154 ? pht_4_122 : _GEN_1209; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1211 = 3'h4 == pht_rindex & 7'h7b == _GEN_9154 ? pht_4_123 : _GEN_1210; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1212 = 3'h4 == pht_rindex & 7'h7c == _GEN_9154 ? pht_4_124 : _GEN_1211; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1213 = 3'h4 == pht_rindex & 7'h7d == _GEN_9154 ? pht_4_125 : _GEN_1212; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1214 = 3'h4 == pht_rindex & 7'h7e == _GEN_9154 ? pht_4_126 : _GEN_1213; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1215 = 3'h4 == pht_rindex & 7'h7f == _GEN_9154 ? pht_4_127 : _GEN_1214; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1216 = 3'h4 == pht_rindex & 8'h80 == _GEN_9346 ? pht_4_128 : _GEN_1215; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1217 = 3'h4 == pht_rindex & 8'h81 == _GEN_9346 ? pht_4_129 : _GEN_1216; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1218 = 3'h4 == pht_rindex & 8'h82 == _GEN_9346 ? pht_4_130 : _GEN_1217; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1219 = 3'h4 == pht_rindex & 8'h83 == _GEN_9346 ? pht_4_131 : _GEN_1218; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1220 = 3'h4 == pht_rindex & 8'h84 == _GEN_9346 ? pht_4_132 : _GEN_1219; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1221 = 3'h4 == pht_rindex & 8'h85 == _GEN_9346 ? pht_4_133 : _GEN_1220; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1222 = 3'h4 == pht_rindex & 8'h86 == _GEN_9346 ? pht_4_134 : _GEN_1221; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1223 = 3'h4 == pht_rindex & 8'h87 == _GEN_9346 ? pht_4_135 : _GEN_1222; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1224 = 3'h4 == pht_rindex & 8'h88 == _GEN_9346 ? pht_4_136 : _GEN_1223; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1225 = 3'h4 == pht_rindex & 8'h89 == _GEN_9346 ? pht_4_137 : _GEN_1224; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1226 = 3'h4 == pht_rindex & 8'h8a == _GEN_9346 ? pht_4_138 : _GEN_1225; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1227 = 3'h4 == pht_rindex & 8'h8b == _GEN_9346 ? pht_4_139 : _GEN_1226; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1228 = 3'h4 == pht_rindex & 8'h8c == _GEN_9346 ? pht_4_140 : _GEN_1227; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1229 = 3'h4 == pht_rindex & 8'h8d == _GEN_9346 ? pht_4_141 : _GEN_1228; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1230 = 3'h4 == pht_rindex & 8'h8e == _GEN_9346 ? pht_4_142 : _GEN_1229; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1231 = 3'h4 == pht_rindex & 8'h8f == _GEN_9346 ? pht_4_143 : _GEN_1230; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1232 = 3'h4 == pht_rindex & 8'h90 == _GEN_9346 ? pht_4_144 : _GEN_1231; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1233 = 3'h4 == pht_rindex & 8'h91 == _GEN_9346 ? pht_4_145 : _GEN_1232; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1234 = 3'h4 == pht_rindex & 8'h92 == _GEN_9346 ? pht_4_146 : _GEN_1233; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1235 = 3'h4 == pht_rindex & 8'h93 == _GEN_9346 ? pht_4_147 : _GEN_1234; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1236 = 3'h4 == pht_rindex & 8'h94 == _GEN_9346 ? pht_4_148 : _GEN_1235; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1237 = 3'h4 == pht_rindex & 8'h95 == _GEN_9346 ? pht_4_149 : _GEN_1236; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1238 = 3'h4 == pht_rindex & 8'h96 == _GEN_9346 ? pht_4_150 : _GEN_1237; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1239 = 3'h4 == pht_rindex & 8'h97 == _GEN_9346 ? pht_4_151 : _GEN_1238; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1240 = 3'h4 == pht_rindex & 8'h98 == _GEN_9346 ? pht_4_152 : _GEN_1239; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1241 = 3'h4 == pht_rindex & 8'h99 == _GEN_9346 ? pht_4_153 : _GEN_1240; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1242 = 3'h4 == pht_rindex & 8'h9a == _GEN_9346 ? pht_4_154 : _GEN_1241; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1243 = 3'h4 == pht_rindex & 8'h9b == _GEN_9346 ? pht_4_155 : _GEN_1242; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1244 = 3'h4 == pht_rindex & 8'h9c == _GEN_9346 ? pht_4_156 : _GEN_1243; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1245 = 3'h4 == pht_rindex & 8'h9d == _GEN_9346 ? pht_4_157 : _GEN_1244; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1246 = 3'h4 == pht_rindex & 8'h9e == _GEN_9346 ? pht_4_158 : _GEN_1245; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1247 = 3'h4 == pht_rindex & 8'h9f == _GEN_9346 ? pht_4_159 : _GEN_1246; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1248 = 3'h4 == pht_rindex & 8'ha0 == _GEN_9346 ? pht_4_160 : _GEN_1247; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1249 = 3'h4 == pht_rindex & 8'ha1 == _GEN_9346 ? pht_4_161 : _GEN_1248; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1250 = 3'h4 == pht_rindex & 8'ha2 == _GEN_9346 ? pht_4_162 : _GEN_1249; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1251 = 3'h4 == pht_rindex & 8'ha3 == _GEN_9346 ? pht_4_163 : _GEN_1250; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1252 = 3'h4 == pht_rindex & 8'ha4 == _GEN_9346 ? pht_4_164 : _GEN_1251; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1253 = 3'h4 == pht_rindex & 8'ha5 == _GEN_9346 ? pht_4_165 : _GEN_1252; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1254 = 3'h4 == pht_rindex & 8'ha6 == _GEN_9346 ? pht_4_166 : _GEN_1253; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1255 = 3'h4 == pht_rindex & 8'ha7 == _GEN_9346 ? pht_4_167 : _GEN_1254; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1256 = 3'h4 == pht_rindex & 8'ha8 == _GEN_9346 ? pht_4_168 : _GEN_1255; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1257 = 3'h4 == pht_rindex & 8'ha9 == _GEN_9346 ? pht_4_169 : _GEN_1256; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1258 = 3'h4 == pht_rindex & 8'haa == _GEN_9346 ? pht_4_170 : _GEN_1257; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1259 = 3'h4 == pht_rindex & 8'hab == _GEN_9346 ? pht_4_171 : _GEN_1258; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1260 = 3'h4 == pht_rindex & 8'hac == _GEN_9346 ? pht_4_172 : _GEN_1259; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1261 = 3'h4 == pht_rindex & 8'had == _GEN_9346 ? pht_4_173 : _GEN_1260; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1262 = 3'h4 == pht_rindex & 8'hae == _GEN_9346 ? pht_4_174 : _GEN_1261; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1263 = 3'h4 == pht_rindex & 8'haf == _GEN_9346 ? pht_4_175 : _GEN_1262; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1264 = 3'h4 == pht_rindex & 8'hb0 == _GEN_9346 ? pht_4_176 : _GEN_1263; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1265 = 3'h4 == pht_rindex & 8'hb1 == _GEN_9346 ? pht_4_177 : _GEN_1264; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1266 = 3'h4 == pht_rindex & 8'hb2 == _GEN_9346 ? pht_4_178 : _GEN_1265; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1267 = 3'h4 == pht_rindex & 8'hb3 == _GEN_9346 ? pht_4_179 : _GEN_1266; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1268 = 3'h4 == pht_rindex & 8'hb4 == _GEN_9346 ? pht_4_180 : _GEN_1267; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1269 = 3'h4 == pht_rindex & 8'hb5 == _GEN_9346 ? pht_4_181 : _GEN_1268; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1270 = 3'h4 == pht_rindex & 8'hb6 == _GEN_9346 ? pht_4_182 : _GEN_1269; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1271 = 3'h4 == pht_rindex & 8'hb7 == _GEN_9346 ? pht_4_183 : _GEN_1270; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1272 = 3'h4 == pht_rindex & 8'hb8 == _GEN_9346 ? pht_4_184 : _GEN_1271; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1273 = 3'h4 == pht_rindex & 8'hb9 == _GEN_9346 ? pht_4_185 : _GEN_1272; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1274 = 3'h4 == pht_rindex & 8'hba == _GEN_9346 ? pht_4_186 : _GEN_1273; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1275 = 3'h4 == pht_rindex & 8'hbb == _GEN_9346 ? pht_4_187 : _GEN_1274; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1276 = 3'h4 == pht_rindex & 8'hbc == _GEN_9346 ? pht_4_188 : _GEN_1275; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1277 = 3'h4 == pht_rindex & 8'hbd == _GEN_9346 ? pht_4_189 : _GEN_1276; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1278 = 3'h4 == pht_rindex & 8'hbe == _GEN_9346 ? pht_4_190 : _GEN_1277; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1279 = 3'h4 == pht_rindex & 8'hbf == _GEN_9346 ? pht_4_191 : _GEN_1278; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1280 = 3'h4 == pht_rindex & 8'hc0 == _GEN_9346 ? pht_4_192 : _GEN_1279; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1281 = 3'h4 == pht_rindex & 8'hc1 == _GEN_9346 ? pht_4_193 : _GEN_1280; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1282 = 3'h4 == pht_rindex & 8'hc2 == _GEN_9346 ? pht_4_194 : _GEN_1281; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1283 = 3'h4 == pht_rindex & 8'hc3 == _GEN_9346 ? pht_4_195 : _GEN_1282; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1284 = 3'h4 == pht_rindex & 8'hc4 == _GEN_9346 ? pht_4_196 : _GEN_1283; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1285 = 3'h4 == pht_rindex & 8'hc5 == _GEN_9346 ? pht_4_197 : _GEN_1284; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1286 = 3'h4 == pht_rindex & 8'hc6 == _GEN_9346 ? pht_4_198 : _GEN_1285; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1287 = 3'h4 == pht_rindex & 8'hc7 == _GEN_9346 ? pht_4_199 : _GEN_1286; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1288 = 3'h4 == pht_rindex & 8'hc8 == _GEN_9346 ? pht_4_200 : _GEN_1287; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1289 = 3'h4 == pht_rindex & 8'hc9 == _GEN_9346 ? pht_4_201 : _GEN_1288; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1290 = 3'h4 == pht_rindex & 8'hca == _GEN_9346 ? pht_4_202 : _GEN_1289; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1291 = 3'h4 == pht_rindex & 8'hcb == _GEN_9346 ? pht_4_203 : _GEN_1290; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1292 = 3'h4 == pht_rindex & 8'hcc == _GEN_9346 ? pht_4_204 : _GEN_1291; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1293 = 3'h4 == pht_rindex & 8'hcd == _GEN_9346 ? pht_4_205 : _GEN_1292; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1294 = 3'h4 == pht_rindex & 8'hce == _GEN_9346 ? pht_4_206 : _GEN_1293; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1295 = 3'h4 == pht_rindex & 8'hcf == _GEN_9346 ? pht_4_207 : _GEN_1294; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1296 = 3'h4 == pht_rindex & 8'hd0 == _GEN_9346 ? pht_4_208 : _GEN_1295; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1297 = 3'h4 == pht_rindex & 8'hd1 == _GEN_9346 ? pht_4_209 : _GEN_1296; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1298 = 3'h4 == pht_rindex & 8'hd2 == _GEN_9346 ? pht_4_210 : _GEN_1297; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1299 = 3'h4 == pht_rindex & 8'hd3 == _GEN_9346 ? pht_4_211 : _GEN_1298; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1300 = 3'h4 == pht_rindex & 8'hd4 == _GEN_9346 ? pht_4_212 : _GEN_1299; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1301 = 3'h4 == pht_rindex & 8'hd5 == _GEN_9346 ? pht_4_213 : _GEN_1300; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1302 = 3'h4 == pht_rindex & 8'hd6 == _GEN_9346 ? pht_4_214 : _GEN_1301; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1303 = 3'h4 == pht_rindex & 8'hd7 == _GEN_9346 ? pht_4_215 : _GEN_1302; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1304 = 3'h4 == pht_rindex & 8'hd8 == _GEN_9346 ? pht_4_216 : _GEN_1303; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1305 = 3'h4 == pht_rindex & 8'hd9 == _GEN_9346 ? pht_4_217 : _GEN_1304; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1306 = 3'h4 == pht_rindex & 8'hda == _GEN_9346 ? pht_4_218 : _GEN_1305; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1307 = 3'h4 == pht_rindex & 8'hdb == _GEN_9346 ? pht_4_219 : _GEN_1306; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1308 = 3'h4 == pht_rindex & 8'hdc == _GEN_9346 ? pht_4_220 : _GEN_1307; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1309 = 3'h4 == pht_rindex & 8'hdd == _GEN_9346 ? pht_4_221 : _GEN_1308; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1310 = 3'h4 == pht_rindex & 8'hde == _GEN_9346 ? pht_4_222 : _GEN_1309; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1311 = 3'h4 == pht_rindex & 8'hdf == _GEN_9346 ? pht_4_223 : _GEN_1310; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1312 = 3'h4 == pht_rindex & 8'he0 == _GEN_9346 ? pht_4_224 : _GEN_1311; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1313 = 3'h4 == pht_rindex & 8'he1 == _GEN_9346 ? pht_4_225 : _GEN_1312; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1314 = 3'h4 == pht_rindex & 8'he2 == _GEN_9346 ? pht_4_226 : _GEN_1313; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1315 = 3'h4 == pht_rindex & 8'he3 == _GEN_9346 ? pht_4_227 : _GEN_1314; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1316 = 3'h4 == pht_rindex & 8'he4 == _GEN_9346 ? pht_4_228 : _GEN_1315; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1317 = 3'h4 == pht_rindex & 8'he5 == _GEN_9346 ? pht_4_229 : _GEN_1316; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1318 = 3'h4 == pht_rindex & 8'he6 == _GEN_9346 ? pht_4_230 : _GEN_1317; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1319 = 3'h4 == pht_rindex & 8'he7 == _GEN_9346 ? pht_4_231 : _GEN_1318; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1320 = 3'h4 == pht_rindex & 8'he8 == _GEN_9346 ? pht_4_232 : _GEN_1319; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1321 = 3'h4 == pht_rindex & 8'he9 == _GEN_9346 ? pht_4_233 : _GEN_1320; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1322 = 3'h4 == pht_rindex & 8'hea == _GEN_9346 ? pht_4_234 : _GEN_1321; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1323 = 3'h4 == pht_rindex & 8'heb == _GEN_9346 ? pht_4_235 : _GEN_1322; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1324 = 3'h4 == pht_rindex & 8'hec == _GEN_9346 ? pht_4_236 : _GEN_1323; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1325 = 3'h4 == pht_rindex & 8'hed == _GEN_9346 ? pht_4_237 : _GEN_1324; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1326 = 3'h4 == pht_rindex & 8'hee == _GEN_9346 ? pht_4_238 : _GEN_1325; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1327 = 3'h4 == pht_rindex & 8'hef == _GEN_9346 ? pht_4_239 : _GEN_1326; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1328 = 3'h4 == pht_rindex & 8'hf0 == _GEN_9346 ? pht_4_240 : _GEN_1327; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1329 = 3'h4 == pht_rindex & 8'hf1 == _GEN_9346 ? pht_4_241 : _GEN_1328; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1330 = 3'h4 == pht_rindex & 8'hf2 == _GEN_9346 ? pht_4_242 : _GEN_1329; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1331 = 3'h4 == pht_rindex & 8'hf3 == _GEN_9346 ? pht_4_243 : _GEN_1330; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1332 = 3'h4 == pht_rindex & 8'hf4 == _GEN_9346 ? pht_4_244 : _GEN_1331; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1333 = 3'h4 == pht_rindex & 8'hf5 == _GEN_9346 ? pht_4_245 : _GEN_1332; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1334 = 3'h4 == pht_rindex & 8'hf6 == _GEN_9346 ? pht_4_246 : _GEN_1333; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1335 = 3'h4 == pht_rindex & 8'hf7 == _GEN_9346 ? pht_4_247 : _GEN_1334; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1336 = 3'h4 == pht_rindex & 8'hf8 == _GEN_9346 ? pht_4_248 : _GEN_1335; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1337 = 3'h4 == pht_rindex & 8'hf9 == _GEN_9346 ? pht_4_249 : _GEN_1336; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1338 = 3'h4 == pht_rindex & 8'hfa == _GEN_9346 ? pht_4_250 : _GEN_1337; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1339 = 3'h4 == pht_rindex & 8'hfb == _GEN_9346 ? pht_4_251 : _GEN_1338; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1340 = 3'h4 == pht_rindex & 8'hfc == _GEN_9346 ? pht_4_252 : _GEN_1339; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1341 = 3'h4 == pht_rindex & 8'hfd == _GEN_9346 ? pht_4_253 : _GEN_1340; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1342 = 3'h4 == pht_rindex & 8'hfe == _GEN_9346 ? pht_4_254 : _GEN_1341; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1343 = 3'h4 == pht_rindex & 8'hff == _GEN_9346 ? pht_4_255 : _GEN_1342; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1344 = 3'h5 == pht_rindex & 6'h0 == pht_raddr ? pht_5_0 : _GEN_1343; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1345 = 3'h5 == pht_rindex & 6'h1 == pht_raddr ? pht_5_1 : _GEN_1344; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1346 = 3'h5 == pht_rindex & 6'h2 == pht_raddr ? pht_5_2 : _GEN_1345; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1347 = 3'h5 == pht_rindex & 6'h3 == pht_raddr ? pht_5_3 : _GEN_1346; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1348 = 3'h5 == pht_rindex & 6'h4 == pht_raddr ? pht_5_4 : _GEN_1347; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1349 = 3'h5 == pht_rindex & 6'h5 == pht_raddr ? pht_5_5 : _GEN_1348; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1350 = 3'h5 == pht_rindex & 6'h6 == pht_raddr ? pht_5_6 : _GEN_1349; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1351 = 3'h5 == pht_rindex & 6'h7 == pht_raddr ? pht_5_7 : _GEN_1350; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1352 = 3'h5 == pht_rindex & 6'h8 == pht_raddr ? pht_5_8 : _GEN_1351; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1353 = 3'h5 == pht_rindex & 6'h9 == pht_raddr ? pht_5_9 : _GEN_1352; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1354 = 3'h5 == pht_rindex & 6'ha == pht_raddr ? pht_5_10 : _GEN_1353; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1355 = 3'h5 == pht_rindex & 6'hb == pht_raddr ? pht_5_11 : _GEN_1354; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1356 = 3'h5 == pht_rindex & 6'hc == pht_raddr ? pht_5_12 : _GEN_1355; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1357 = 3'h5 == pht_rindex & 6'hd == pht_raddr ? pht_5_13 : _GEN_1356; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1358 = 3'h5 == pht_rindex & 6'he == pht_raddr ? pht_5_14 : _GEN_1357; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1359 = 3'h5 == pht_rindex & 6'hf == pht_raddr ? pht_5_15 : _GEN_1358; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1360 = 3'h5 == pht_rindex & 6'h10 == pht_raddr ? pht_5_16 : _GEN_1359; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1361 = 3'h5 == pht_rindex & 6'h11 == pht_raddr ? pht_5_17 : _GEN_1360; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1362 = 3'h5 == pht_rindex & 6'h12 == pht_raddr ? pht_5_18 : _GEN_1361; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1363 = 3'h5 == pht_rindex & 6'h13 == pht_raddr ? pht_5_19 : _GEN_1362; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1364 = 3'h5 == pht_rindex & 6'h14 == pht_raddr ? pht_5_20 : _GEN_1363; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1365 = 3'h5 == pht_rindex & 6'h15 == pht_raddr ? pht_5_21 : _GEN_1364; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1366 = 3'h5 == pht_rindex & 6'h16 == pht_raddr ? pht_5_22 : _GEN_1365; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1367 = 3'h5 == pht_rindex & 6'h17 == pht_raddr ? pht_5_23 : _GEN_1366; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1368 = 3'h5 == pht_rindex & 6'h18 == pht_raddr ? pht_5_24 : _GEN_1367; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1369 = 3'h5 == pht_rindex & 6'h19 == pht_raddr ? pht_5_25 : _GEN_1368; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1370 = 3'h5 == pht_rindex & 6'h1a == pht_raddr ? pht_5_26 : _GEN_1369; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1371 = 3'h5 == pht_rindex & 6'h1b == pht_raddr ? pht_5_27 : _GEN_1370; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1372 = 3'h5 == pht_rindex & 6'h1c == pht_raddr ? pht_5_28 : _GEN_1371; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1373 = 3'h5 == pht_rindex & 6'h1d == pht_raddr ? pht_5_29 : _GEN_1372; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1374 = 3'h5 == pht_rindex & 6'h1e == pht_raddr ? pht_5_30 : _GEN_1373; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1375 = 3'h5 == pht_rindex & 6'h1f == pht_raddr ? pht_5_31 : _GEN_1374; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1376 = 3'h5 == pht_rindex & 6'h20 == pht_raddr ? pht_5_32 : _GEN_1375; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1377 = 3'h5 == pht_rindex & 6'h21 == pht_raddr ? pht_5_33 : _GEN_1376; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1378 = 3'h5 == pht_rindex & 6'h22 == pht_raddr ? pht_5_34 : _GEN_1377; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1379 = 3'h5 == pht_rindex & 6'h23 == pht_raddr ? pht_5_35 : _GEN_1378; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1380 = 3'h5 == pht_rindex & 6'h24 == pht_raddr ? pht_5_36 : _GEN_1379; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1381 = 3'h5 == pht_rindex & 6'h25 == pht_raddr ? pht_5_37 : _GEN_1380; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1382 = 3'h5 == pht_rindex & 6'h26 == pht_raddr ? pht_5_38 : _GEN_1381; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1383 = 3'h5 == pht_rindex & 6'h27 == pht_raddr ? pht_5_39 : _GEN_1382; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1384 = 3'h5 == pht_rindex & 6'h28 == pht_raddr ? pht_5_40 : _GEN_1383; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1385 = 3'h5 == pht_rindex & 6'h29 == pht_raddr ? pht_5_41 : _GEN_1384; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1386 = 3'h5 == pht_rindex & 6'h2a == pht_raddr ? pht_5_42 : _GEN_1385; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1387 = 3'h5 == pht_rindex & 6'h2b == pht_raddr ? pht_5_43 : _GEN_1386; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1388 = 3'h5 == pht_rindex & 6'h2c == pht_raddr ? pht_5_44 : _GEN_1387; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1389 = 3'h5 == pht_rindex & 6'h2d == pht_raddr ? pht_5_45 : _GEN_1388; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1390 = 3'h5 == pht_rindex & 6'h2e == pht_raddr ? pht_5_46 : _GEN_1389; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1391 = 3'h5 == pht_rindex & 6'h2f == pht_raddr ? pht_5_47 : _GEN_1390; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1392 = 3'h5 == pht_rindex & 6'h30 == pht_raddr ? pht_5_48 : _GEN_1391; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1393 = 3'h5 == pht_rindex & 6'h31 == pht_raddr ? pht_5_49 : _GEN_1392; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1394 = 3'h5 == pht_rindex & 6'h32 == pht_raddr ? pht_5_50 : _GEN_1393; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1395 = 3'h5 == pht_rindex & 6'h33 == pht_raddr ? pht_5_51 : _GEN_1394; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1396 = 3'h5 == pht_rindex & 6'h34 == pht_raddr ? pht_5_52 : _GEN_1395; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1397 = 3'h5 == pht_rindex & 6'h35 == pht_raddr ? pht_5_53 : _GEN_1396; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1398 = 3'h5 == pht_rindex & 6'h36 == pht_raddr ? pht_5_54 : _GEN_1397; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1399 = 3'h5 == pht_rindex & 6'h37 == pht_raddr ? pht_5_55 : _GEN_1398; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1400 = 3'h5 == pht_rindex & 6'h38 == pht_raddr ? pht_5_56 : _GEN_1399; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1401 = 3'h5 == pht_rindex & 6'h39 == pht_raddr ? pht_5_57 : _GEN_1400; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1402 = 3'h5 == pht_rindex & 6'h3a == pht_raddr ? pht_5_58 : _GEN_1401; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1403 = 3'h5 == pht_rindex & 6'h3b == pht_raddr ? pht_5_59 : _GEN_1402; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1404 = 3'h5 == pht_rindex & 6'h3c == pht_raddr ? pht_5_60 : _GEN_1403; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1405 = 3'h5 == pht_rindex & 6'h3d == pht_raddr ? pht_5_61 : _GEN_1404; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1406 = 3'h5 == pht_rindex & 6'h3e == pht_raddr ? pht_5_62 : _GEN_1405; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1407 = 3'h5 == pht_rindex & 6'h3f == pht_raddr ? pht_5_63 : _GEN_1406; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1408 = 3'h5 == pht_rindex & 7'h40 == _GEN_9154 ? pht_5_64 : _GEN_1407; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1409 = 3'h5 == pht_rindex & 7'h41 == _GEN_9154 ? pht_5_65 : _GEN_1408; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1410 = 3'h5 == pht_rindex & 7'h42 == _GEN_9154 ? pht_5_66 : _GEN_1409; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1411 = 3'h5 == pht_rindex & 7'h43 == _GEN_9154 ? pht_5_67 : _GEN_1410; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1412 = 3'h5 == pht_rindex & 7'h44 == _GEN_9154 ? pht_5_68 : _GEN_1411; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1413 = 3'h5 == pht_rindex & 7'h45 == _GEN_9154 ? pht_5_69 : _GEN_1412; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1414 = 3'h5 == pht_rindex & 7'h46 == _GEN_9154 ? pht_5_70 : _GEN_1413; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1415 = 3'h5 == pht_rindex & 7'h47 == _GEN_9154 ? pht_5_71 : _GEN_1414; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1416 = 3'h5 == pht_rindex & 7'h48 == _GEN_9154 ? pht_5_72 : _GEN_1415; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1417 = 3'h5 == pht_rindex & 7'h49 == _GEN_9154 ? pht_5_73 : _GEN_1416; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1418 = 3'h5 == pht_rindex & 7'h4a == _GEN_9154 ? pht_5_74 : _GEN_1417; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1419 = 3'h5 == pht_rindex & 7'h4b == _GEN_9154 ? pht_5_75 : _GEN_1418; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1420 = 3'h5 == pht_rindex & 7'h4c == _GEN_9154 ? pht_5_76 : _GEN_1419; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1421 = 3'h5 == pht_rindex & 7'h4d == _GEN_9154 ? pht_5_77 : _GEN_1420; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1422 = 3'h5 == pht_rindex & 7'h4e == _GEN_9154 ? pht_5_78 : _GEN_1421; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1423 = 3'h5 == pht_rindex & 7'h4f == _GEN_9154 ? pht_5_79 : _GEN_1422; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1424 = 3'h5 == pht_rindex & 7'h50 == _GEN_9154 ? pht_5_80 : _GEN_1423; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1425 = 3'h5 == pht_rindex & 7'h51 == _GEN_9154 ? pht_5_81 : _GEN_1424; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1426 = 3'h5 == pht_rindex & 7'h52 == _GEN_9154 ? pht_5_82 : _GEN_1425; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1427 = 3'h5 == pht_rindex & 7'h53 == _GEN_9154 ? pht_5_83 : _GEN_1426; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1428 = 3'h5 == pht_rindex & 7'h54 == _GEN_9154 ? pht_5_84 : _GEN_1427; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1429 = 3'h5 == pht_rindex & 7'h55 == _GEN_9154 ? pht_5_85 : _GEN_1428; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1430 = 3'h5 == pht_rindex & 7'h56 == _GEN_9154 ? pht_5_86 : _GEN_1429; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1431 = 3'h5 == pht_rindex & 7'h57 == _GEN_9154 ? pht_5_87 : _GEN_1430; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1432 = 3'h5 == pht_rindex & 7'h58 == _GEN_9154 ? pht_5_88 : _GEN_1431; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1433 = 3'h5 == pht_rindex & 7'h59 == _GEN_9154 ? pht_5_89 : _GEN_1432; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1434 = 3'h5 == pht_rindex & 7'h5a == _GEN_9154 ? pht_5_90 : _GEN_1433; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1435 = 3'h5 == pht_rindex & 7'h5b == _GEN_9154 ? pht_5_91 : _GEN_1434; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1436 = 3'h5 == pht_rindex & 7'h5c == _GEN_9154 ? pht_5_92 : _GEN_1435; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1437 = 3'h5 == pht_rindex & 7'h5d == _GEN_9154 ? pht_5_93 : _GEN_1436; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1438 = 3'h5 == pht_rindex & 7'h5e == _GEN_9154 ? pht_5_94 : _GEN_1437; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1439 = 3'h5 == pht_rindex & 7'h5f == _GEN_9154 ? pht_5_95 : _GEN_1438; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1440 = 3'h5 == pht_rindex & 7'h60 == _GEN_9154 ? pht_5_96 : _GEN_1439; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1441 = 3'h5 == pht_rindex & 7'h61 == _GEN_9154 ? pht_5_97 : _GEN_1440; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1442 = 3'h5 == pht_rindex & 7'h62 == _GEN_9154 ? pht_5_98 : _GEN_1441; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1443 = 3'h5 == pht_rindex & 7'h63 == _GEN_9154 ? pht_5_99 : _GEN_1442; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1444 = 3'h5 == pht_rindex & 7'h64 == _GEN_9154 ? pht_5_100 : _GEN_1443; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1445 = 3'h5 == pht_rindex & 7'h65 == _GEN_9154 ? pht_5_101 : _GEN_1444; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1446 = 3'h5 == pht_rindex & 7'h66 == _GEN_9154 ? pht_5_102 : _GEN_1445; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1447 = 3'h5 == pht_rindex & 7'h67 == _GEN_9154 ? pht_5_103 : _GEN_1446; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1448 = 3'h5 == pht_rindex & 7'h68 == _GEN_9154 ? pht_5_104 : _GEN_1447; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1449 = 3'h5 == pht_rindex & 7'h69 == _GEN_9154 ? pht_5_105 : _GEN_1448; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1450 = 3'h5 == pht_rindex & 7'h6a == _GEN_9154 ? pht_5_106 : _GEN_1449; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1451 = 3'h5 == pht_rindex & 7'h6b == _GEN_9154 ? pht_5_107 : _GEN_1450; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1452 = 3'h5 == pht_rindex & 7'h6c == _GEN_9154 ? pht_5_108 : _GEN_1451; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1453 = 3'h5 == pht_rindex & 7'h6d == _GEN_9154 ? pht_5_109 : _GEN_1452; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1454 = 3'h5 == pht_rindex & 7'h6e == _GEN_9154 ? pht_5_110 : _GEN_1453; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1455 = 3'h5 == pht_rindex & 7'h6f == _GEN_9154 ? pht_5_111 : _GEN_1454; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1456 = 3'h5 == pht_rindex & 7'h70 == _GEN_9154 ? pht_5_112 : _GEN_1455; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1457 = 3'h5 == pht_rindex & 7'h71 == _GEN_9154 ? pht_5_113 : _GEN_1456; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1458 = 3'h5 == pht_rindex & 7'h72 == _GEN_9154 ? pht_5_114 : _GEN_1457; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1459 = 3'h5 == pht_rindex & 7'h73 == _GEN_9154 ? pht_5_115 : _GEN_1458; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1460 = 3'h5 == pht_rindex & 7'h74 == _GEN_9154 ? pht_5_116 : _GEN_1459; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1461 = 3'h5 == pht_rindex & 7'h75 == _GEN_9154 ? pht_5_117 : _GEN_1460; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1462 = 3'h5 == pht_rindex & 7'h76 == _GEN_9154 ? pht_5_118 : _GEN_1461; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1463 = 3'h5 == pht_rindex & 7'h77 == _GEN_9154 ? pht_5_119 : _GEN_1462; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1464 = 3'h5 == pht_rindex & 7'h78 == _GEN_9154 ? pht_5_120 : _GEN_1463; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1465 = 3'h5 == pht_rindex & 7'h79 == _GEN_9154 ? pht_5_121 : _GEN_1464; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1466 = 3'h5 == pht_rindex & 7'h7a == _GEN_9154 ? pht_5_122 : _GEN_1465; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1467 = 3'h5 == pht_rindex & 7'h7b == _GEN_9154 ? pht_5_123 : _GEN_1466; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1468 = 3'h5 == pht_rindex & 7'h7c == _GEN_9154 ? pht_5_124 : _GEN_1467; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1469 = 3'h5 == pht_rindex & 7'h7d == _GEN_9154 ? pht_5_125 : _GEN_1468; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1470 = 3'h5 == pht_rindex & 7'h7e == _GEN_9154 ? pht_5_126 : _GEN_1469; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1471 = 3'h5 == pht_rindex & 7'h7f == _GEN_9154 ? pht_5_127 : _GEN_1470; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1472 = 3'h5 == pht_rindex & 8'h80 == _GEN_9346 ? pht_5_128 : _GEN_1471; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1473 = 3'h5 == pht_rindex & 8'h81 == _GEN_9346 ? pht_5_129 : _GEN_1472; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1474 = 3'h5 == pht_rindex & 8'h82 == _GEN_9346 ? pht_5_130 : _GEN_1473; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1475 = 3'h5 == pht_rindex & 8'h83 == _GEN_9346 ? pht_5_131 : _GEN_1474; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1476 = 3'h5 == pht_rindex & 8'h84 == _GEN_9346 ? pht_5_132 : _GEN_1475; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1477 = 3'h5 == pht_rindex & 8'h85 == _GEN_9346 ? pht_5_133 : _GEN_1476; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1478 = 3'h5 == pht_rindex & 8'h86 == _GEN_9346 ? pht_5_134 : _GEN_1477; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1479 = 3'h5 == pht_rindex & 8'h87 == _GEN_9346 ? pht_5_135 : _GEN_1478; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1480 = 3'h5 == pht_rindex & 8'h88 == _GEN_9346 ? pht_5_136 : _GEN_1479; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1481 = 3'h5 == pht_rindex & 8'h89 == _GEN_9346 ? pht_5_137 : _GEN_1480; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1482 = 3'h5 == pht_rindex & 8'h8a == _GEN_9346 ? pht_5_138 : _GEN_1481; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1483 = 3'h5 == pht_rindex & 8'h8b == _GEN_9346 ? pht_5_139 : _GEN_1482; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1484 = 3'h5 == pht_rindex & 8'h8c == _GEN_9346 ? pht_5_140 : _GEN_1483; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1485 = 3'h5 == pht_rindex & 8'h8d == _GEN_9346 ? pht_5_141 : _GEN_1484; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1486 = 3'h5 == pht_rindex & 8'h8e == _GEN_9346 ? pht_5_142 : _GEN_1485; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1487 = 3'h5 == pht_rindex & 8'h8f == _GEN_9346 ? pht_5_143 : _GEN_1486; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1488 = 3'h5 == pht_rindex & 8'h90 == _GEN_9346 ? pht_5_144 : _GEN_1487; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1489 = 3'h5 == pht_rindex & 8'h91 == _GEN_9346 ? pht_5_145 : _GEN_1488; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1490 = 3'h5 == pht_rindex & 8'h92 == _GEN_9346 ? pht_5_146 : _GEN_1489; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1491 = 3'h5 == pht_rindex & 8'h93 == _GEN_9346 ? pht_5_147 : _GEN_1490; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1492 = 3'h5 == pht_rindex & 8'h94 == _GEN_9346 ? pht_5_148 : _GEN_1491; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1493 = 3'h5 == pht_rindex & 8'h95 == _GEN_9346 ? pht_5_149 : _GEN_1492; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1494 = 3'h5 == pht_rindex & 8'h96 == _GEN_9346 ? pht_5_150 : _GEN_1493; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1495 = 3'h5 == pht_rindex & 8'h97 == _GEN_9346 ? pht_5_151 : _GEN_1494; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1496 = 3'h5 == pht_rindex & 8'h98 == _GEN_9346 ? pht_5_152 : _GEN_1495; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1497 = 3'h5 == pht_rindex & 8'h99 == _GEN_9346 ? pht_5_153 : _GEN_1496; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1498 = 3'h5 == pht_rindex & 8'h9a == _GEN_9346 ? pht_5_154 : _GEN_1497; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1499 = 3'h5 == pht_rindex & 8'h9b == _GEN_9346 ? pht_5_155 : _GEN_1498; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1500 = 3'h5 == pht_rindex & 8'h9c == _GEN_9346 ? pht_5_156 : _GEN_1499; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1501 = 3'h5 == pht_rindex & 8'h9d == _GEN_9346 ? pht_5_157 : _GEN_1500; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1502 = 3'h5 == pht_rindex & 8'h9e == _GEN_9346 ? pht_5_158 : _GEN_1501; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1503 = 3'h5 == pht_rindex & 8'h9f == _GEN_9346 ? pht_5_159 : _GEN_1502; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1504 = 3'h5 == pht_rindex & 8'ha0 == _GEN_9346 ? pht_5_160 : _GEN_1503; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1505 = 3'h5 == pht_rindex & 8'ha1 == _GEN_9346 ? pht_5_161 : _GEN_1504; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1506 = 3'h5 == pht_rindex & 8'ha2 == _GEN_9346 ? pht_5_162 : _GEN_1505; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1507 = 3'h5 == pht_rindex & 8'ha3 == _GEN_9346 ? pht_5_163 : _GEN_1506; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1508 = 3'h5 == pht_rindex & 8'ha4 == _GEN_9346 ? pht_5_164 : _GEN_1507; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1509 = 3'h5 == pht_rindex & 8'ha5 == _GEN_9346 ? pht_5_165 : _GEN_1508; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1510 = 3'h5 == pht_rindex & 8'ha6 == _GEN_9346 ? pht_5_166 : _GEN_1509; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1511 = 3'h5 == pht_rindex & 8'ha7 == _GEN_9346 ? pht_5_167 : _GEN_1510; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1512 = 3'h5 == pht_rindex & 8'ha8 == _GEN_9346 ? pht_5_168 : _GEN_1511; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1513 = 3'h5 == pht_rindex & 8'ha9 == _GEN_9346 ? pht_5_169 : _GEN_1512; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1514 = 3'h5 == pht_rindex & 8'haa == _GEN_9346 ? pht_5_170 : _GEN_1513; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1515 = 3'h5 == pht_rindex & 8'hab == _GEN_9346 ? pht_5_171 : _GEN_1514; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1516 = 3'h5 == pht_rindex & 8'hac == _GEN_9346 ? pht_5_172 : _GEN_1515; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1517 = 3'h5 == pht_rindex & 8'had == _GEN_9346 ? pht_5_173 : _GEN_1516; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1518 = 3'h5 == pht_rindex & 8'hae == _GEN_9346 ? pht_5_174 : _GEN_1517; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1519 = 3'h5 == pht_rindex & 8'haf == _GEN_9346 ? pht_5_175 : _GEN_1518; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1520 = 3'h5 == pht_rindex & 8'hb0 == _GEN_9346 ? pht_5_176 : _GEN_1519; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1521 = 3'h5 == pht_rindex & 8'hb1 == _GEN_9346 ? pht_5_177 : _GEN_1520; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1522 = 3'h5 == pht_rindex & 8'hb2 == _GEN_9346 ? pht_5_178 : _GEN_1521; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1523 = 3'h5 == pht_rindex & 8'hb3 == _GEN_9346 ? pht_5_179 : _GEN_1522; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1524 = 3'h5 == pht_rindex & 8'hb4 == _GEN_9346 ? pht_5_180 : _GEN_1523; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1525 = 3'h5 == pht_rindex & 8'hb5 == _GEN_9346 ? pht_5_181 : _GEN_1524; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1526 = 3'h5 == pht_rindex & 8'hb6 == _GEN_9346 ? pht_5_182 : _GEN_1525; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1527 = 3'h5 == pht_rindex & 8'hb7 == _GEN_9346 ? pht_5_183 : _GEN_1526; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1528 = 3'h5 == pht_rindex & 8'hb8 == _GEN_9346 ? pht_5_184 : _GEN_1527; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1529 = 3'h5 == pht_rindex & 8'hb9 == _GEN_9346 ? pht_5_185 : _GEN_1528; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1530 = 3'h5 == pht_rindex & 8'hba == _GEN_9346 ? pht_5_186 : _GEN_1529; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1531 = 3'h5 == pht_rindex & 8'hbb == _GEN_9346 ? pht_5_187 : _GEN_1530; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1532 = 3'h5 == pht_rindex & 8'hbc == _GEN_9346 ? pht_5_188 : _GEN_1531; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1533 = 3'h5 == pht_rindex & 8'hbd == _GEN_9346 ? pht_5_189 : _GEN_1532; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1534 = 3'h5 == pht_rindex & 8'hbe == _GEN_9346 ? pht_5_190 : _GEN_1533; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1535 = 3'h5 == pht_rindex & 8'hbf == _GEN_9346 ? pht_5_191 : _GEN_1534; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1536 = 3'h5 == pht_rindex & 8'hc0 == _GEN_9346 ? pht_5_192 : _GEN_1535; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1537 = 3'h5 == pht_rindex & 8'hc1 == _GEN_9346 ? pht_5_193 : _GEN_1536; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1538 = 3'h5 == pht_rindex & 8'hc2 == _GEN_9346 ? pht_5_194 : _GEN_1537; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1539 = 3'h5 == pht_rindex & 8'hc3 == _GEN_9346 ? pht_5_195 : _GEN_1538; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1540 = 3'h5 == pht_rindex & 8'hc4 == _GEN_9346 ? pht_5_196 : _GEN_1539; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1541 = 3'h5 == pht_rindex & 8'hc5 == _GEN_9346 ? pht_5_197 : _GEN_1540; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1542 = 3'h5 == pht_rindex & 8'hc6 == _GEN_9346 ? pht_5_198 : _GEN_1541; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1543 = 3'h5 == pht_rindex & 8'hc7 == _GEN_9346 ? pht_5_199 : _GEN_1542; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1544 = 3'h5 == pht_rindex & 8'hc8 == _GEN_9346 ? pht_5_200 : _GEN_1543; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1545 = 3'h5 == pht_rindex & 8'hc9 == _GEN_9346 ? pht_5_201 : _GEN_1544; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1546 = 3'h5 == pht_rindex & 8'hca == _GEN_9346 ? pht_5_202 : _GEN_1545; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1547 = 3'h5 == pht_rindex & 8'hcb == _GEN_9346 ? pht_5_203 : _GEN_1546; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1548 = 3'h5 == pht_rindex & 8'hcc == _GEN_9346 ? pht_5_204 : _GEN_1547; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1549 = 3'h5 == pht_rindex & 8'hcd == _GEN_9346 ? pht_5_205 : _GEN_1548; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1550 = 3'h5 == pht_rindex & 8'hce == _GEN_9346 ? pht_5_206 : _GEN_1549; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1551 = 3'h5 == pht_rindex & 8'hcf == _GEN_9346 ? pht_5_207 : _GEN_1550; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1552 = 3'h5 == pht_rindex & 8'hd0 == _GEN_9346 ? pht_5_208 : _GEN_1551; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1553 = 3'h5 == pht_rindex & 8'hd1 == _GEN_9346 ? pht_5_209 : _GEN_1552; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1554 = 3'h5 == pht_rindex & 8'hd2 == _GEN_9346 ? pht_5_210 : _GEN_1553; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1555 = 3'h5 == pht_rindex & 8'hd3 == _GEN_9346 ? pht_5_211 : _GEN_1554; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1556 = 3'h5 == pht_rindex & 8'hd4 == _GEN_9346 ? pht_5_212 : _GEN_1555; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1557 = 3'h5 == pht_rindex & 8'hd5 == _GEN_9346 ? pht_5_213 : _GEN_1556; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1558 = 3'h5 == pht_rindex & 8'hd6 == _GEN_9346 ? pht_5_214 : _GEN_1557; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1559 = 3'h5 == pht_rindex & 8'hd7 == _GEN_9346 ? pht_5_215 : _GEN_1558; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1560 = 3'h5 == pht_rindex & 8'hd8 == _GEN_9346 ? pht_5_216 : _GEN_1559; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1561 = 3'h5 == pht_rindex & 8'hd9 == _GEN_9346 ? pht_5_217 : _GEN_1560; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1562 = 3'h5 == pht_rindex & 8'hda == _GEN_9346 ? pht_5_218 : _GEN_1561; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1563 = 3'h5 == pht_rindex & 8'hdb == _GEN_9346 ? pht_5_219 : _GEN_1562; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1564 = 3'h5 == pht_rindex & 8'hdc == _GEN_9346 ? pht_5_220 : _GEN_1563; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1565 = 3'h5 == pht_rindex & 8'hdd == _GEN_9346 ? pht_5_221 : _GEN_1564; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1566 = 3'h5 == pht_rindex & 8'hde == _GEN_9346 ? pht_5_222 : _GEN_1565; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1567 = 3'h5 == pht_rindex & 8'hdf == _GEN_9346 ? pht_5_223 : _GEN_1566; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1568 = 3'h5 == pht_rindex & 8'he0 == _GEN_9346 ? pht_5_224 : _GEN_1567; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1569 = 3'h5 == pht_rindex & 8'he1 == _GEN_9346 ? pht_5_225 : _GEN_1568; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1570 = 3'h5 == pht_rindex & 8'he2 == _GEN_9346 ? pht_5_226 : _GEN_1569; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1571 = 3'h5 == pht_rindex & 8'he3 == _GEN_9346 ? pht_5_227 : _GEN_1570; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1572 = 3'h5 == pht_rindex & 8'he4 == _GEN_9346 ? pht_5_228 : _GEN_1571; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1573 = 3'h5 == pht_rindex & 8'he5 == _GEN_9346 ? pht_5_229 : _GEN_1572; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1574 = 3'h5 == pht_rindex & 8'he6 == _GEN_9346 ? pht_5_230 : _GEN_1573; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1575 = 3'h5 == pht_rindex & 8'he7 == _GEN_9346 ? pht_5_231 : _GEN_1574; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1576 = 3'h5 == pht_rindex & 8'he8 == _GEN_9346 ? pht_5_232 : _GEN_1575; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1577 = 3'h5 == pht_rindex & 8'he9 == _GEN_9346 ? pht_5_233 : _GEN_1576; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1578 = 3'h5 == pht_rindex & 8'hea == _GEN_9346 ? pht_5_234 : _GEN_1577; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1579 = 3'h5 == pht_rindex & 8'heb == _GEN_9346 ? pht_5_235 : _GEN_1578; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1580 = 3'h5 == pht_rindex & 8'hec == _GEN_9346 ? pht_5_236 : _GEN_1579; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1581 = 3'h5 == pht_rindex & 8'hed == _GEN_9346 ? pht_5_237 : _GEN_1580; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1582 = 3'h5 == pht_rindex & 8'hee == _GEN_9346 ? pht_5_238 : _GEN_1581; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1583 = 3'h5 == pht_rindex & 8'hef == _GEN_9346 ? pht_5_239 : _GEN_1582; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1584 = 3'h5 == pht_rindex & 8'hf0 == _GEN_9346 ? pht_5_240 : _GEN_1583; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1585 = 3'h5 == pht_rindex & 8'hf1 == _GEN_9346 ? pht_5_241 : _GEN_1584; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1586 = 3'h5 == pht_rindex & 8'hf2 == _GEN_9346 ? pht_5_242 : _GEN_1585; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1587 = 3'h5 == pht_rindex & 8'hf3 == _GEN_9346 ? pht_5_243 : _GEN_1586; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1588 = 3'h5 == pht_rindex & 8'hf4 == _GEN_9346 ? pht_5_244 : _GEN_1587; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1589 = 3'h5 == pht_rindex & 8'hf5 == _GEN_9346 ? pht_5_245 : _GEN_1588; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1590 = 3'h5 == pht_rindex & 8'hf6 == _GEN_9346 ? pht_5_246 : _GEN_1589; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1591 = 3'h5 == pht_rindex & 8'hf7 == _GEN_9346 ? pht_5_247 : _GEN_1590; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1592 = 3'h5 == pht_rindex & 8'hf8 == _GEN_9346 ? pht_5_248 : _GEN_1591; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1593 = 3'h5 == pht_rindex & 8'hf9 == _GEN_9346 ? pht_5_249 : _GEN_1592; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1594 = 3'h5 == pht_rindex & 8'hfa == _GEN_9346 ? pht_5_250 : _GEN_1593; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1595 = 3'h5 == pht_rindex & 8'hfb == _GEN_9346 ? pht_5_251 : _GEN_1594; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1596 = 3'h5 == pht_rindex & 8'hfc == _GEN_9346 ? pht_5_252 : _GEN_1595; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1597 = 3'h5 == pht_rindex & 8'hfd == _GEN_9346 ? pht_5_253 : _GEN_1596; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1598 = 3'h5 == pht_rindex & 8'hfe == _GEN_9346 ? pht_5_254 : _GEN_1597; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1599 = 3'h5 == pht_rindex & 8'hff == _GEN_9346 ? pht_5_255 : _GEN_1598; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1600 = 3'h6 == pht_rindex & 6'h0 == pht_raddr ? pht_6_0 : _GEN_1599; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1601 = 3'h6 == pht_rindex & 6'h1 == pht_raddr ? pht_6_1 : _GEN_1600; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1602 = 3'h6 == pht_rindex & 6'h2 == pht_raddr ? pht_6_2 : _GEN_1601; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1603 = 3'h6 == pht_rindex & 6'h3 == pht_raddr ? pht_6_3 : _GEN_1602; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1604 = 3'h6 == pht_rindex & 6'h4 == pht_raddr ? pht_6_4 : _GEN_1603; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1605 = 3'h6 == pht_rindex & 6'h5 == pht_raddr ? pht_6_5 : _GEN_1604; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1606 = 3'h6 == pht_rindex & 6'h6 == pht_raddr ? pht_6_6 : _GEN_1605; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1607 = 3'h6 == pht_rindex & 6'h7 == pht_raddr ? pht_6_7 : _GEN_1606; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1608 = 3'h6 == pht_rindex & 6'h8 == pht_raddr ? pht_6_8 : _GEN_1607; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1609 = 3'h6 == pht_rindex & 6'h9 == pht_raddr ? pht_6_9 : _GEN_1608; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1610 = 3'h6 == pht_rindex & 6'ha == pht_raddr ? pht_6_10 : _GEN_1609; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1611 = 3'h6 == pht_rindex & 6'hb == pht_raddr ? pht_6_11 : _GEN_1610; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1612 = 3'h6 == pht_rindex & 6'hc == pht_raddr ? pht_6_12 : _GEN_1611; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1613 = 3'h6 == pht_rindex & 6'hd == pht_raddr ? pht_6_13 : _GEN_1612; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1614 = 3'h6 == pht_rindex & 6'he == pht_raddr ? pht_6_14 : _GEN_1613; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1615 = 3'h6 == pht_rindex & 6'hf == pht_raddr ? pht_6_15 : _GEN_1614; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1616 = 3'h6 == pht_rindex & 6'h10 == pht_raddr ? pht_6_16 : _GEN_1615; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1617 = 3'h6 == pht_rindex & 6'h11 == pht_raddr ? pht_6_17 : _GEN_1616; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1618 = 3'h6 == pht_rindex & 6'h12 == pht_raddr ? pht_6_18 : _GEN_1617; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1619 = 3'h6 == pht_rindex & 6'h13 == pht_raddr ? pht_6_19 : _GEN_1618; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1620 = 3'h6 == pht_rindex & 6'h14 == pht_raddr ? pht_6_20 : _GEN_1619; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1621 = 3'h6 == pht_rindex & 6'h15 == pht_raddr ? pht_6_21 : _GEN_1620; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1622 = 3'h6 == pht_rindex & 6'h16 == pht_raddr ? pht_6_22 : _GEN_1621; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1623 = 3'h6 == pht_rindex & 6'h17 == pht_raddr ? pht_6_23 : _GEN_1622; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1624 = 3'h6 == pht_rindex & 6'h18 == pht_raddr ? pht_6_24 : _GEN_1623; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1625 = 3'h6 == pht_rindex & 6'h19 == pht_raddr ? pht_6_25 : _GEN_1624; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1626 = 3'h6 == pht_rindex & 6'h1a == pht_raddr ? pht_6_26 : _GEN_1625; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1627 = 3'h6 == pht_rindex & 6'h1b == pht_raddr ? pht_6_27 : _GEN_1626; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1628 = 3'h6 == pht_rindex & 6'h1c == pht_raddr ? pht_6_28 : _GEN_1627; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1629 = 3'h6 == pht_rindex & 6'h1d == pht_raddr ? pht_6_29 : _GEN_1628; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1630 = 3'h6 == pht_rindex & 6'h1e == pht_raddr ? pht_6_30 : _GEN_1629; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1631 = 3'h6 == pht_rindex & 6'h1f == pht_raddr ? pht_6_31 : _GEN_1630; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1632 = 3'h6 == pht_rindex & 6'h20 == pht_raddr ? pht_6_32 : _GEN_1631; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1633 = 3'h6 == pht_rindex & 6'h21 == pht_raddr ? pht_6_33 : _GEN_1632; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1634 = 3'h6 == pht_rindex & 6'h22 == pht_raddr ? pht_6_34 : _GEN_1633; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1635 = 3'h6 == pht_rindex & 6'h23 == pht_raddr ? pht_6_35 : _GEN_1634; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1636 = 3'h6 == pht_rindex & 6'h24 == pht_raddr ? pht_6_36 : _GEN_1635; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1637 = 3'h6 == pht_rindex & 6'h25 == pht_raddr ? pht_6_37 : _GEN_1636; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1638 = 3'h6 == pht_rindex & 6'h26 == pht_raddr ? pht_6_38 : _GEN_1637; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1639 = 3'h6 == pht_rindex & 6'h27 == pht_raddr ? pht_6_39 : _GEN_1638; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1640 = 3'h6 == pht_rindex & 6'h28 == pht_raddr ? pht_6_40 : _GEN_1639; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1641 = 3'h6 == pht_rindex & 6'h29 == pht_raddr ? pht_6_41 : _GEN_1640; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1642 = 3'h6 == pht_rindex & 6'h2a == pht_raddr ? pht_6_42 : _GEN_1641; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1643 = 3'h6 == pht_rindex & 6'h2b == pht_raddr ? pht_6_43 : _GEN_1642; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1644 = 3'h6 == pht_rindex & 6'h2c == pht_raddr ? pht_6_44 : _GEN_1643; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1645 = 3'h6 == pht_rindex & 6'h2d == pht_raddr ? pht_6_45 : _GEN_1644; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1646 = 3'h6 == pht_rindex & 6'h2e == pht_raddr ? pht_6_46 : _GEN_1645; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1647 = 3'h6 == pht_rindex & 6'h2f == pht_raddr ? pht_6_47 : _GEN_1646; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1648 = 3'h6 == pht_rindex & 6'h30 == pht_raddr ? pht_6_48 : _GEN_1647; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1649 = 3'h6 == pht_rindex & 6'h31 == pht_raddr ? pht_6_49 : _GEN_1648; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1650 = 3'h6 == pht_rindex & 6'h32 == pht_raddr ? pht_6_50 : _GEN_1649; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1651 = 3'h6 == pht_rindex & 6'h33 == pht_raddr ? pht_6_51 : _GEN_1650; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1652 = 3'h6 == pht_rindex & 6'h34 == pht_raddr ? pht_6_52 : _GEN_1651; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1653 = 3'h6 == pht_rindex & 6'h35 == pht_raddr ? pht_6_53 : _GEN_1652; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1654 = 3'h6 == pht_rindex & 6'h36 == pht_raddr ? pht_6_54 : _GEN_1653; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1655 = 3'h6 == pht_rindex & 6'h37 == pht_raddr ? pht_6_55 : _GEN_1654; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1656 = 3'h6 == pht_rindex & 6'h38 == pht_raddr ? pht_6_56 : _GEN_1655; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1657 = 3'h6 == pht_rindex & 6'h39 == pht_raddr ? pht_6_57 : _GEN_1656; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1658 = 3'h6 == pht_rindex & 6'h3a == pht_raddr ? pht_6_58 : _GEN_1657; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1659 = 3'h6 == pht_rindex & 6'h3b == pht_raddr ? pht_6_59 : _GEN_1658; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1660 = 3'h6 == pht_rindex & 6'h3c == pht_raddr ? pht_6_60 : _GEN_1659; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1661 = 3'h6 == pht_rindex & 6'h3d == pht_raddr ? pht_6_61 : _GEN_1660; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1662 = 3'h6 == pht_rindex & 6'h3e == pht_raddr ? pht_6_62 : _GEN_1661; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1663 = 3'h6 == pht_rindex & 6'h3f == pht_raddr ? pht_6_63 : _GEN_1662; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1664 = 3'h6 == pht_rindex & 7'h40 == _GEN_9154 ? pht_6_64 : _GEN_1663; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1665 = 3'h6 == pht_rindex & 7'h41 == _GEN_9154 ? pht_6_65 : _GEN_1664; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1666 = 3'h6 == pht_rindex & 7'h42 == _GEN_9154 ? pht_6_66 : _GEN_1665; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1667 = 3'h6 == pht_rindex & 7'h43 == _GEN_9154 ? pht_6_67 : _GEN_1666; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1668 = 3'h6 == pht_rindex & 7'h44 == _GEN_9154 ? pht_6_68 : _GEN_1667; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1669 = 3'h6 == pht_rindex & 7'h45 == _GEN_9154 ? pht_6_69 : _GEN_1668; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1670 = 3'h6 == pht_rindex & 7'h46 == _GEN_9154 ? pht_6_70 : _GEN_1669; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1671 = 3'h6 == pht_rindex & 7'h47 == _GEN_9154 ? pht_6_71 : _GEN_1670; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1672 = 3'h6 == pht_rindex & 7'h48 == _GEN_9154 ? pht_6_72 : _GEN_1671; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1673 = 3'h6 == pht_rindex & 7'h49 == _GEN_9154 ? pht_6_73 : _GEN_1672; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1674 = 3'h6 == pht_rindex & 7'h4a == _GEN_9154 ? pht_6_74 : _GEN_1673; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1675 = 3'h6 == pht_rindex & 7'h4b == _GEN_9154 ? pht_6_75 : _GEN_1674; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1676 = 3'h6 == pht_rindex & 7'h4c == _GEN_9154 ? pht_6_76 : _GEN_1675; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1677 = 3'h6 == pht_rindex & 7'h4d == _GEN_9154 ? pht_6_77 : _GEN_1676; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1678 = 3'h6 == pht_rindex & 7'h4e == _GEN_9154 ? pht_6_78 : _GEN_1677; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1679 = 3'h6 == pht_rindex & 7'h4f == _GEN_9154 ? pht_6_79 : _GEN_1678; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1680 = 3'h6 == pht_rindex & 7'h50 == _GEN_9154 ? pht_6_80 : _GEN_1679; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1681 = 3'h6 == pht_rindex & 7'h51 == _GEN_9154 ? pht_6_81 : _GEN_1680; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1682 = 3'h6 == pht_rindex & 7'h52 == _GEN_9154 ? pht_6_82 : _GEN_1681; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1683 = 3'h6 == pht_rindex & 7'h53 == _GEN_9154 ? pht_6_83 : _GEN_1682; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1684 = 3'h6 == pht_rindex & 7'h54 == _GEN_9154 ? pht_6_84 : _GEN_1683; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1685 = 3'h6 == pht_rindex & 7'h55 == _GEN_9154 ? pht_6_85 : _GEN_1684; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1686 = 3'h6 == pht_rindex & 7'h56 == _GEN_9154 ? pht_6_86 : _GEN_1685; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1687 = 3'h6 == pht_rindex & 7'h57 == _GEN_9154 ? pht_6_87 : _GEN_1686; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1688 = 3'h6 == pht_rindex & 7'h58 == _GEN_9154 ? pht_6_88 : _GEN_1687; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1689 = 3'h6 == pht_rindex & 7'h59 == _GEN_9154 ? pht_6_89 : _GEN_1688; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1690 = 3'h6 == pht_rindex & 7'h5a == _GEN_9154 ? pht_6_90 : _GEN_1689; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1691 = 3'h6 == pht_rindex & 7'h5b == _GEN_9154 ? pht_6_91 : _GEN_1690; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1692 = 3'h6 == pht_rindex & 7'h5c == _GEN_9154 ? pht_6_92 : _GEN_1691; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1693 = 3'h6 == pht_rindex & 7'h5d == _GEN_9154 ? pht_6_93 : _GEN_1692; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1694 = 3'h6 == pht_rindex & 7'h5e == _GEN_9154 ? pht_6_94 : _GEN_1693; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1695 = 3'h6 == pht_rindex & 7'h5f == _GEN_9154 ? pht_6_95 : _GEN_1694; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1696 = 3'h6 == pht_rindex & 7'h60 == _GEN_9154 ? pht_6_96 : _GEN_1695; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1697 = 3'h6 == pht_rindex & 7'h61 == _GEN_9154 ? pht_6_97 : _GEN_1696; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1698 = 3'h6 == pht_rindex & 7'h62 == _GEN_9154 ? pht_6_98 : _GEN_1697; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1699 = 3'h6 == pht_rindex & 7'h63 == _GEN_9154 ? pht_6_99 : _GEN_1698; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1700 = 3'h6 == pht_rindex & 7'h64 == _GEN_9154 ? pht_6_100 : _GEN_1699; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1701 = 3'h6 == pht_rindex & 7'h65 == _GEN_9154 ? pht_6_101 : _GEN_1700; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1702 = 3'h6 == pht_rindex & 7'h66 == _GEN_9154 ? pht_6_102 : _GEN_1701; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1703 = 3'h6 == pht_rindex & 7'h67 == _GEN_9154 ? pht_6_103 : _GEN_1702; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1704 = 3'h6 == pht_rindex & 7'h68 == _GEN_9154 ? pht_6_104 : _GEN_1703; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1705 = 3'h6 == pht_rindex & 7'h69 == _GEN_9154 ? pht_6_105 : _GEN_1704; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1706 = 3'h6 == pht_rindex & 7'h6a == _GEN_9154 ? pht_6_106 : _GEN_1705; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1707 = 3'h6 == pht_rindex & 7'h6b == _GEN_9154 ? pht_6_107 : _GEN_1706; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1708 = 3'h6 == pht_rindex & 7'h6c == _GEN_9154 ? pht_6_108 : _GEN_1707; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1709 = 3'h6 == pht_rindex & 7'h6d == _GEN_9154 ? pht_6_109 : _GEN_1708; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1710 = 3'h6 == pht_rindex & 7'h6e == _GEN_9154 ? pht_6_110 : _GEN_1709; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1711 = 3'h6 == pht_rindex & 7'h6f == _GEN_9154 ? pht_6_111 : _GEN_1710; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1712 = 3'h6 == pht_rindex & 7'h70 == _GEN_9154 ? pht_6_112 : _GEN_1711; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1713 = 3'h6 == pht_rindex & 7'h71 == _GEN_9154 ? pht_6_113 : _GEN_1712; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1714 = 3'h6 == pht_rindex & 7'h72 == _GEN_9154 ? pht_6_114 : _GEN_1713; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1715 = 3'h6 == pht_rindex & 7'h73 == _GEN_9154 ? pht_6_115 : _GEN_1714; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1716 = 3'h6 == pht_rindex & 7'h74 == _GEN_9154 ? pht_6_116 : _GEN_1715; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1717 = 3'h6 == pht_rindex & 7'h75 == _GEN_9154 ? pht_6_117 : _GEN_1716; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1718 = 3'h6 == pht_rindex & 7'h76 == _GEN_9154 ? pht_6_118 : _GEN_1717; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1719 = 3'h6 == pht_rindex & 7'h77 == _GEN_9154 ? pht_6_119 : _GEN_1718; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1720 = 3'h6 == pht_rindex & 7'h78 == _GEN_9154 ? pht_6_120 : _GEN_1719; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1721 = 3'h6 == pht_rindex & 7'h79 == _GEN_9154 ? pht_6_121 : _GEN_1720; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1722 = 3'h6 == pht_rindex & 7'h7a == _GEN_9154 ? pht_6_122 : _GEN_1721; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1723 = 3'h6 == pht_rindex & 7'h7b == _GEN_9154 ? pht_6_123 : _GEN_1722; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1724 = 3'h6 == pht_rindex & 7'h7c == _GEN_9154 ? pht_6_124 : _GEN_1723; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1725 = 3'h6 == pht_rindex & 7'h7d == _GEN_9154 ? pht_6_125 : _GEN_1724; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1726 = 3'h6 == pht_rindex & 7'h7e == _GEN_9154 ? pht_6_126 : _GEN_1725; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1727 = 3'h6 == pht_rindex & 7'h7f == _GEN_9154 ? pht_6_127 : _GEN_1726; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1728 = 3'h6 == pht_rindex & 8'h80 == _GEN_9346 ? pht_6_128 : _GEN_1727; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1729 = 3'h6 == pht_rindex & 8'h81 == _GEN_9346 ? pht_6_129 : _GEN_1728; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1730 = 3'h6 == pht_rindex & 8'h82 == _GEN_9346 ? pht_6_130 : _GEN_1729; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1731 = 3'h6 == pht_rindex & 8'h83 == _GEN_9346 ? pht_6_131 : _GEN_1730; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1732 = 3'h6 == pht_rindex & 8'h84 == _GEN_9346 ? pht_6_132 : _GEN_1731; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1733 = 3'h6 == pht_rindex & 8'h85 == _GEN_9346 ? pht_6_133 : _GEN_1732; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1734 = 3'h6 == pht_rindex & 8'h86 == _GEN_9346 ? pht_6_134 : _GEN_1733; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1735 = 3'h6 == pht_rindex & 8'h87 == _GEN_9346 ? pht_6_135 : _GEN_1734; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1736 = 3'h6 == pht_rindex & 8'h88 == _GEN_9346 ? pht_6_136 : _GEN_1735; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1737 = 3'h6 == pht_rindex & 8'h89 == _GEN_9346 ? pht_6_137 : _GEN_1736; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1738 = 3'h6 == pht_rindex & 8'h8a == _GEN_9346 ? pht_6_138 : _GEN_1737; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1739 = 3'h6 == pht_rindex & 8'h8b == _GEN_9346 ? pht_6_139 : _GEN_1738; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1740 = 3'h6 == pht_rindex & 8'h8c == _GEN_9346 ? pht_6_140 : _GEN_1739; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1741 = 3'h6 == pht_rindex & 8'h8d == _GEN_9346 ? pht_6_141 : _GEN_1740; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1742 = 3'h6 == pht_rindex & 8'h8e == _GEN_9346 ? pht_6_142 : _GEN_1741; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1743 = 3'h6 == pht_rindex & 8'h8f == _GEN_9346 ? pht_6_143 : _GEN_1742; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1744 = 3'h6 == pht_rindex & 8'h90 == _GEN_9346 ? pht_6_144 : _GEN_1743; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1745 = 3'h6 == pht_rindex & 8'h91 == _GEN_9346 ? pht_6_145 : _GEN_1744; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1746 = 3'h6 == pht_rindex & 8'h92 == _GEN_9346 ? pht_6_146 : _GEN_1745; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1747 = 3'h6 == pht_rindex & 8'h93 == _GEN_9346 ? pht_6_147 : _GEN_1746; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1748 = 3'h6 == pht_rindex & 8'h94 == _GEN_9346 ? pht_6_148 : _GEN_1747; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1749 = 3'h6 == pht_rindex & 8'h95 == _GEN_9346 ? pht_6_149 : _GEN_1748; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1750 = 3'h6 == pht_rindex & 8'h96 == _GEN_9346 ? pht_6_150 : _GEN_1749; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1751 = 3'h6 == pht_rindex & 8'h97 == _GEN_9346 ? pht_6_151 : _GEN_1750; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1752 = 3'h6 == pht_rindex & 8'h98 == _GEN_9346 ? pht_6_152 : _GEN_1751; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1753 = 3'h6 == pht_rindex & 8'h99 == _GEN_9346 ? pht_6_153 : _GEN_1752; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1754 = 3'h6 == pht_rindex & 8'h9a == _GEN_9346 ? pht_6_154 : _GEN_1753; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1755 = 3'h6 == pht_rindex & 8'h9b == _GEN_9346 ? pht_6_155 : _GEN_1754; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1756 = 3'h6 == pht_rindex & 8'h9c == _GEN_9346 ? pht_6_156 : _GEN_1755; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1757 = 3'h6 == pht_rindex & 8'h9d == _GEN_9346 ? pht_6_157 : _GEN_1756; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1758 = 3'h6 == pht_rindex & 8'h9e == _GEN_9346 ? pht_6_158 : _GEN_1757; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1759 = 3'h6 == pht_rindex & 8'h9f == _GEN_9346 ? pht_6_159 : _GEN_1758; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1760 = 3'h6 == pht_rindex & 8'ha0 == _GEN_9346 ? pht_6_160 : _GEN_1759; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1761 = 3'h6 == pht_rindex & 8'ha1 == _GEN_9346 ? pht_6_161 : _GEN_1760; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1762 = 3'h6 == pht_rindex & 8'ha2 == _GEN_9346 ? pht_6_162 : _GEN_1761; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1763 = 3'h6 == pht_rindex & 8'ha3 == _GEN_9346 ? pht_6_163 : _GEN_1762; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1764 = 3'h6 == pht_rindex & 8'ha4 == _GEN_9346 ? pht_6_164 : _GEN_1763; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1765 = 3'h6 == pht_rindex & 8'ha5 == _GEN_9346 ? pht_6_165 : _GEN_1764; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1766 = 3'h6 == pht_rindex & 8'ha6 == _GEN_9346 ? pht_6_166 : _GEN_1765; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1767 = 3'h6 == pht_rindex & 8'ha7 == _GEN_9346 ? pht_6_167 : _GEN_1766; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1768 = 3'h6 == pht_rindex & 8'ha8 == _GEN_9346 ? pht_6_168 : _GEN_1767; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1769 = 3'h6 == pht_rindex & 8'ha9 == _GEN_9346 ? pht_6_169 : _GEN_1768; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1770 = 3'h6 == pht_rindex & 8'haa == _GEN_9346 ? pht_6_170 : _GEN_1769; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1771 = 3'h6 == pht_rindex & 8'hab == _GEN_9346 ? pht_6_171 : _GEN_1770; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1772 = 3'h6 == pht_rindex & 8'hac == _GEN_9346 ? pht_6_172 : _GEN_1771; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1773 = 3'h6 == pht_rindex & 8'had == _GEN_9346 ? pht_6_173 : _GEN_1772; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1774 = 3'h6 == pht_rindex & 8'hae == _GEN_9346 ? pht_6_174 : _GEN_1773; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1775 = 3'h6 == pht_rindex & 8'haf == _GEN_9346 ? pht_6_175 : _GEN_1774; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1776 = 3'h6 == pht_rindex & 8'hb0 == _GEN_9346 ? pht_6_176 : _GEN_1775; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1777 = 3'h6 == pht_rindex & 8'hb1 == _GEN_9346 ? pht_6_177 : _GEN_1776; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1778 = 3'h6 == pht_rindex & 8'hb2 == _GEN_9346 ? pht_6_178 : _GEN_1777; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1779 = 3'h6 == pht_rindex & 8'hb3 == _GEN_9346 ? pht_6_179 : _GEN_1778; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1780 = 3'h6 == pht_rindex & 8'hb4 == _GEN_9346 ? pht_6_180 : _GEN_1779; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1781 = 3'h6 == pht_rindex & 8'hb5 == _GEN_9346 ? pht_6_181 : _GEN_1780; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1782 = 3'h6 == pht_rindex & 8'hb6 == _GEN_9346 ? pht_6_182 : _GEN_1781; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1783 = 3'h6 == pht_rindex & 8'hb7 == _GEN_9346 ? pht_6_183 : _GEN_1782; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1784 = 3'h6 == pht_rindex & 8'hb8 == _GEN_9346 ? pht_6_184 : _GEN_1783; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1785 = 3'h6 == pht_rindex & 8'hb9 == _GEN_9346 ? pht_6_185 : _GEN_1784; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1786 = 3'h6 == pht_rindex & 8'hba == _GEN_9346 ? pht_6_186 : _GEN_1785; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1787 = 3'h6 == pht_rindex & 8'hbb == _GEN_9346 ? pht_6_187 : _GEN_1786; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1788 = 3'h6 == pht_rindex & 8'hbc == _GEN_9346 ? pht_6_188 : _GEN_1787; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1789 = 3'h6 == pht_rindex & 8'hbd == _GEN_9346 ? pht_6_189 : _GEN_1788; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1790 = 3'h6 == pht_rindex & 8'hbe == _GEN_9346 ? pht_6_190 : _GEN_1789; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1791 = 3'h6 == pht_rindex & 8'hbf == _GEN_9346 ? pht_6_191 : _GEN_1790; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1792 = 3'h6 == pht_rindex & 8'hc0 == _GEN_9346 ? pht_6_192 : _GEN_1791; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1793 = 3'h6 == pht_rindex & 8'hc1 == _GEN_9346 ? pht_6_193 : _GEN_1792; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1794 = 3'h6 == pht_rindex & 8'hc2 == _GEN_9346 ? pht_6_194 : _GEN_1793; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1795 = 3'h6 == pht_rindex & 8'hc3 == _GEN_9346 ? pht_6_195 : _GEN_1794; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1796 = 3'h6 == pht_rindex & 8'hc4 == _GEN_9346 ? pht_6_196 : _GEN_1795; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1797 = 3'h6 == pht_rindex & 8'hc5 == _GEN_9346 ? pht_6_197 : _GEN_1796; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1798 = 3'h6 == pht_rindex & 8'hc6 == _GEN_9346 ? pht_6_198 : _GEN_1797; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1799 = 3'h6 == pht_rindex & 8'hc7 == _GEN_9346 ? pht_6_199 : _GEN_1798; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1800 = 3'h6 == pht_rindex & 8'hc8 == _GEN_9346 ? pht_6_200 : _GEN_1799; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1801 = 3'h6 == pht_rindex & 8'hc9 == _GEN_9346 ? pht_6_201 : _GEN_1800; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1802 = 3'h6 == pht_rindex & 8'hca == _GEN_9346 ? pht_6_202 : _GEN_1801; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1803 = 3'h6 == pht_rindex & 8'hcb == _GEN_9346 ? pht_6_203 : _GEN_1802; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1804 = 3'h6 == pht_rindex & 8'hcc == _GEN_9346 ? pht_6_204 : _GEN_1803; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1805 = 3'h6 == pht_rindex & 8'hcd == _GEN_9346 ? pht_6_205 : _GEN_1804; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1806 = 3'h6 == pht_rindex & 8'hce == _GEN_9346 ? pht_6_206 : _GEN_1805; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1807 = 3'h6 == pht_rindex & 8'hcf == _GEN_9346 ? pht_6_207 : _GEN_1806; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1808 = 3'h6 == pht_rindex & 8'hd0 == _GEN_9346 ? pht_6_208 : _GEN_1807; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1809 = 3'h6 == pht_rindex & 8'hd1 == _GEN_9346 ? pht_6_209 : _GEN_1808; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1810 = 3'h6 == pht_rindex & 8'hd2 == _GEN_9346 ? pht_6_210 : _GEN_1809; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1811 = 3'h6 == pht_rindex & 8'hd3 == _GEN_9346 ? pht_6_211 : _GEN_1810; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1812 = 3'h6 == pht_rindex & 8'hd4 == _GEN_9346 ? pht_6_212 : _GEN_1811; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1813 = 3'h6 == pht_rindex & 8'hd5 == _GEN_9346 ? pht_6_213 : _GEN_1812; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1814 = 3'h6 == pht_rindex & 8'hd6 == _GEN_9346 ? pht_6_214 : _GEN_1813; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1815 = 3'h6 == pht_rindex & 8'hd7 == _GEN_9346 ? pht_6_215 : _GEN_1814; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1816 = 3'h6 == pht_rindex & 8'hd8 == _GEN_9346 ? pht_6_216 : _GEN_1815; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1817 = 3'h6 == pht_rindex & 8'hd9 == _GEN_9346 ? pht_6_217 : _GEN_1816; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1818 = 3'h6 == pht_rindex & 8'hda == _GEN_9346 ? pht_6_218 : _GEN_1817; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1819 = 3'h6 == pht_rindex & 8'hdb == _GEN_9346 ? pht_6_219 : _GEN_1818; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1820 = 3'h6 == pht_rindex & 8'hdc == _GEN_9346 ? pht_6_220 : _GEN_1819; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1821 = 3'h6 == pht_rindex & 8'hdd == _GEN_9346 ? pht_6_221 : _GEN_1820; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1822 = 3'h6 == pht_rindex & 8'hde == _GEN_9346 ? pht_6_222 : _GEN_1821; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1823 = 3'h6 == pht_rindex & 8'hdf == _GEN_9346 ? pht_6_223 : _GEN_1822; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1824 = 3'h6 == pht_rindex & 8'he0 == _GEN_9346 ? pht_6_224 : _GEN_1823; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1825 = 3'h6 == pht_rindex & 8'he1 == _GEN_9346 ? pht_6_225 : _GEN_1824; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1826 = 3'h6 == pht_rindex & 8'he2 == _GEN_9346 ? pht_6_226 : _GEN_1825; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1827 = 3'h6 == pht_rindex & 8'he3 == _GEN_9346 ? pht_6_227 : _GEN_1826; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1828 = 3'h6 == pht_rindex & 8'he4 == _GEN_9346 ? pht_6_228 : _GEN_1827; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1829 = 3'h6 == pht_rindex & 8'he5 == _GEN_9346 ? pht_6_229 : _GEN_1828; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1830 = 3'h6 == pht_rindex & 8'he6 == _GEN_9346 ? pht_6_230 : _GEN_1829; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1831 = 3'h6 == pht_rindex & 8'he7 == _GEN_9346 ? pht_6_231 : _GEN_1830; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1832 = 3'h6 == pht_rindex & 8'he8 == _GEN_9346 ? pht_6_232 : _GEN_1831; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1833 = 3'h6 == pht_rindex & 8'he9 == _GEN_9346 ? pht_6_233 : _GEN_1832; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1834 = 3'h6 == pht_rindex & 8'hea == _GEN_9346 ? pht_6_234 : _GEN_1833; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1835 = 3'h6 == pht_rindex & 8'heb == _GEN_9346 ? pht_6_235 : _GEN_1834; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1836 = 3'h6 == pht_rindex & 8'hec == _GEN_9346 ? pht_6_236 : _GEN_1835; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1837 = 3'h6 == pht_rindex & 8'hed == _GEN_9346 ? pht_6_237 : _GEN_1836; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1838 = 3'h6 == pht_rindex & 8'hee == _GEN_9346 ? pht_6_238 : _GEN_1837; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1839 = 3'h6 == pht_rindex & 8'hef == _GEN_9346 ? pht_6_239 : _GEN_1838; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1840 = 3'h6 == pht_rindex & 8'hf0 == _GEN_9346 ? pht_6_240 : _GEN_1839; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1841 = 3'h6 == pht_rindex & 8'hf1 == _GEN_9346 ? pht_6_241 : _GEN_1840; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1842 = 3'h6 == pht_rindex & 8'hf2 == _GEN_9346 ? pht_6_242 : _GEN_1841; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1843 = 3'h6 == pht_rindex & 8'hf3 == _GEN_9346 ? pht_6_243 : _GEN_1842; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1844 = 3'h6 == pht_rindex & 8'hf4 == _GEN_9346 ? pht_6_244 : _GEN_1843; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1845 = 3'h6 == pht_rindex & 8'hf5 == _GEN_9346 ? pht_6_245 : _GEN_1844; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1846 = 3'h6 == pht_rindex & 8'hf6 == _GEN_9346 ? pht_6_246 : _GEN_1845; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1847 = 3'h6 == pht_rindex & 8'hf7 == _GEN_9346 ? pht_6_247 : _GEN_1846; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1848 = 3'h6 == pht_rindex & 8'hf8 == _GEN_9346 ? pht_6_248 : _GEN_1847; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1849 = 3'h6 == pht_rindex & 8'hf9 == _GEN_9346 ? pht_6_249 : _GEN_1848; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1850 = 3'h6 == pht_rindex & 8'hfa == _GEN_9346 ? pht_6_250 : _GEN_1849; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1851 = 3'h6 == pht_rindex & 8'hfb == _GEN_9346 ? pht_6_251 : _GEN_1850; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1852 = 3'h6 == pht_rindex & 8'hfc == _GEN_9346 ? pht_6_252 : _GEN_1851; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1853 = 3'h6 == pht_rindex & 8'hfd == _GEN_9346 ? pht_6_253 : _GEN_1852; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1854 = 3'h6 == pht_rindex & 8'hfe == _GEN_9346 ? pht_6_254 : _GEN_1853; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1855 = 3'h6 == pht_rindex & 8'hff == _GEN_9346 ? pht_6_255 : _GEN_1854; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1856 = 3'h7 == pht_rindex & 6'h0 == pht_raddr ? pht_7_0 : _GEN_1855; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1857 = 3'h7 == pht_rindex & 6'h1 == pht_raddr ? pht_7_1 : _GEN_1856; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1858 = 3'h7 == pht_rindex & 6'h2 == pht_raddr ? pht_7_2 : _GEN_1857; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1859 = 3'h7 == pht_rindex & 6'h3 == pht_raddr ? pht_7_3 : _GEN_1858; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1860 = 3'h7 == pht_rindex & 6'h4 == pht_raddr ? pht_7_4 : _GEN_1859; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1861 = 3'h7 == pht_rindex & 6'h5 == pht_raddr ? pht_7_5 : _GEN_1860; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1862 = 3'h7 == pht_rindex & 6'h6 == pht_raddr ? pht_7_6 : _GEN_1861; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1863 = 3'h7 == pht_rindex & 6'h7 == pht_raddr ? pht_7_7 : _GEN_1862; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1864 = 3'h7 == pht_rindex & 6'h8 == pht_raddr ? pht_7_8 : _GEN_1863; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1865 = 3'h7 == pht_rindex & 6'h9 == pht_raddr ? pht_7_9 : _GEN_1864; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1866 = 3'h7 == pht_rindex & 6'ha == pht_raddr ? pht_7_10 : _GEN_1865; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1867 = 3'h7 == pht_rindex & 6'hb == pht_raddr ? pht_7_11 : _GEN_1866; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1868 = 3'h7 == pht_rindex & 6'hc == pht_raddr ? pht_7_12 : _GEN_1867; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1869 = 3'h7 == pht_rindex & 6'hd == pht_raddr ? pht_7_13 : _GEN_1868; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1870 = 3'h7 == pht_rindex & 6'he == pht_raddr ? pht_7_14 : _GEN_1869; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1871 = 3'h7 == pht_rindex & 6'hf == pht_raddr ? pht_7_15 : _GEN_1870; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1872 = 3'h7 == pht_rindex & 6'h10 == pht_raddr ? pht_7_16 : _GEN_1871; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1873 = 3'h7 == pht_rindex & 6'h11 == pht_raddr ? pht_7_17 : _GEN_1872; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1874 = 3'h7 == pht_rindex & 6'h12 == pht_raddr ? pht_7_18 : _GEN_1873; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1875 = 3'h7 == pht_rindex & 6'h13 == pht_raddr ? pht_7_19 : _GEN_1874; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1876 = 3'h7 == pht_rindex & 6'h14 == pht_raddr ? pht_7_20 : _GEN_1875; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1877 = 3'h7 == pht_rindex & 6'h15 == pht_raddr ? pht_7_21 : _GEN_1876; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1878 = 3'h7 == pht_rindex & 6'h16 == pht_raddr ? pht_7_22 : _GEN_1877; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1879 = 3'h7 == pht_rindex & 6'h17 == pht_raddr ? pht_7_23 : _GEN_1878; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1880 = 3'h7 == pht_rindex & 6'h18 == pht_raddr ? pht_7_24 : _GEN_1879; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1881 = 3'h7 == pht_rindex & 6'h19 == pht_raddr ? pht_7_25 : _GEN_1880; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1882 = 3'h7 == pht_rindex & 6'h1a == pht_raddr ? pht_7_26 : _GEN_1881; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1883 = 3'h7 == pht_rindex & 6'h1b == pht_raddr ? pht_7_27 : _GEN_1882; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1884 = 3'h7 == pht_rindex & 6'h1c == pht_raddr ? pht_7_28 : _GEN_1883; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1885 = 3'h7 == pht_rindex & 6'h1d == pht_raddr ? pht_7_29 : _GEN_1884; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1886 = 3'h7 == pht_rindex & 6'h1e == pht_raddr ? pht_7_30 : _GEN_1885; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1887 = 3'h7 == pht_rindex & 6'h1f == pht_raddr ? pht_7_31 : _GEN_1886; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1888 = 3'h7 == pht_rindex & 6'h20 == pht_raddr ? pht_7_32 : _GEN_1887; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1889 = 3'h7 == pht_rindex & 6'h21 == pht_raddr ? pht_7_33 : _GEN_1888; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1890 = 3'h7 == pht_rindex & 6'h22 == pht_raddr ? pht_7_34 : _GEN_1889; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1891 = 3'h7 == pht_rindex & 6'h23 == pht_raddr ? pht_7_35 : _GEN_1890; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1892 = 3'h7 == pht_rindex & 6'h24 == pht_raddr ? pht_7_36 : _GEN_1891; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1893 = 3'h7 == pht_rindex & 6'h25 == pht_raddr ? pht_7_37 : _GEN_1892; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1894 = 3'h7 == pht_rindex & 6'h26 == pht_raddr ? pht_7_38 : _GEN_1893; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1895 = 3'h7 == pht_rindex & 6'h27 == pht_raddr ? pht_7_39 : _GEN_1894; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1896 = 3'h7 == pht_rindex & 6'h28 == pht_raddr ? pht_7_40 : _GEN_1895; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1897 = 3'h7 == pht_rindex & 6'h29 == pht_raddr ? pht_7_41 : _GEN_1896; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1898 = 3'h7 == pht_rindex & 6'h2a == pht_raddr ? pht_7_42 : _GEN_1897; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1899 = 3'h7 == pht_rindex & 6'h2b == pht_raddr ? pht_7_43 : _GEN_1898; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1900 = 3'h7 == pht_rindex & 6'h2c == pht_raddr ? pht_7_44 : _GEN_1899; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1901 = 3'h7 == pht_rindex & 6'h2d == pht_raddr ? pht_7_45 : _GEN_1900; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1902 = 3'h7 == pht_rindex & 6'h2e == pht_raddr ? pht_7_46 : _GEN_1901; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1903 = 3'h7 == pht_rindex & 6'h2f == pht_raddr ? pht_7_47 : _GEN_1902; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1904 = 3'h7 == pht_rindex & 6'h30 == pht_raddr ? pht_7_48 : _GEN_1903; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1905 = 3'h7 == pht_rindex & 6'h31 == pht_raddr ? pht_7_49 : _GEN_1904; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1906 = 3'h7 == pht_rindex & 6'h32 == pht_raddr ? pht_7_50 : _GEN_1905; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1907 = 3'h7 == pht_rindex & 6'h33 == pht_raddr ? pht_7_51 : _GEN_1906; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1908 = 3'h7 == pht_rindex & 6'h34 == pht_raddr ? pht_7_52 : _GEN_1907; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1909 = 3'h7 == pht_rindex & 6'h35 == pht_raddr ? pht_7_53 : _GEN_1908; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1910 = 3'h7 == pht_rindex & 6'h36 == pht_raddr ? pht_7_54 : _GEN_1909; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1911 = 3'h7 == pht_rindex & 6'h37 == pht_raddr ? pht_7_55 : _GEN_1910; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1912 = 3'h7 == pht_rindex & 6'h38 == pht_raddr ? pht_7_56 : _GEN_1911; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1913 = 3'h7 == pht_rindex & 6'h39 == pht_raddr ? pht_7_57 : _GEN_1912; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1914 = 3'h7 == pht_rindex & 6'h3a == pht_raddr ? pht_7_58 : _GEN_1913; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1915 = 3'h7 == pht_rindex & 6'h3b == pht_raddr ? pht_7_59 : _GEN_1914; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1916 = 3'h7 == pht_rindex & 6'h3c == pht_raddr ? pht_7_60 : _GEN_1915; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1917 = 3'h7 == pht_rindex & 6'h3d == pht_raddr ? pht_7_61 : _GEN_1916; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1918 = 3'h7 == pht_rindex & 6'h3e == pht_raddr ? pht_7_62 : _GEN_1917; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1919 = 3'h7 == pht_rindex & 6'h3f == pht_raddr ? pht_7_63 : _GEN_1918; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1920 = 3'h7 == pht_rindex & 7'h40 == _GEN_9154 ? pht_7_64 : _GEN_1919; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1921 = 3'h7 == pht_rindex & 7'h41 == _GEN_9154 ? pht_7_65 : _GEN_1920; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1922 = 3'h7 == pht_rindex & 7'h42 == _GEN_9154 ? pht_7_66 : _GEN_1921; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1923 = 3'h7 == pht_rindex & 7'h43 == _GEN_9154 ? pht_7_67 : _GEN_1922; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1924 = 3'h7 == pht_rindex & 7'h44 == _GEN_9154 ? pht_7_68 : _GEN_1923; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1925 = 3'h7 == pht_rindex & 7'h45 == _GEN_9154 ? pht_7_69 : _GEN_1924; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1926 = 3'h7 == pht_rindex & 7'h46 == _GEN_9154 ? pht_7_70 : _GEN_1925; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1927 = 3'h7 == pht_rindex & 7'h47 == _GEN_9154 ? pht_7_71 : _GEN_1926; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1928 = 3'h7 == pht_rindex & 7'h48 == _GEN_9154 ? pht_7_72 : _GEN_1927; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1929 = 3'h7 == pht_rindex & 7'h49 == _GEN_9154 ? pht_7_73 : _GEN_1928; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1930 = 3'h7 == pht_rindex & 7'h4a == _GEN_9154 ? pht_7_74 : _GEN_1929; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1931 = 3'h7 == pht_rindex & 7'h4b == _GEN_9154 ? pht_7_75 : _GEN_1930; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1932 = 3'h7 == pht_rindex & 7'h4c == _GEN_9154 ? pht_7_76 : _GEN_1931; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1933 = 3'h7 == pht_rindex & 7'h4d == _GEN_9154 ? pht_7_77 : _GEN_1932; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1934 = 3'h7 == pht_rindex & 7'h4e == _GEN_9154 ? pht_7_78 : _GEN_1933; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1935 = 3'h7 == pht_rindex & 7'h4f == _GEN_9154 ? pht_7_79 : _GEN_1934; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1936 = 3'h7 == pht_rindex & 7'h50 == _GEN_9154 ? pht_7_80 : _GEN_1935; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1937 = 3'h7 == pht_rindex & 7'h51 == _GEN_9154 ? pht_7_81 : _GEN_1936; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1938 = 3'h7 == pht_rindex & 7'h52 == _GEN_9154 ? pht_7_82 : _GEN_1937; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1939 = 3'h7 == pht_rindex & 7'h53 == _GEN_9154 ? pht_7_83 : _GEN_1938; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1940 = 3'h7 == pht_rindex & 7'h54 == _GEN_9154 ? pht_7_84 : _GEN_1939; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1941 = 3'h7 == pht_rindex & 7'h55 == _GEN_9154 ? pht_7_85 : _GEN_1940; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1942 = 3'h7 == pht_rindex & 7'h56 == _GEN_9154 ? pht_7_86 : _GEN_1941; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1943 = 3'h7 == pht_rindex & 7'h57 == _GEN_9154 ? pht_7_87 : _GEN_1942; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1944 = 3'h7 == pht_rindex & 7'h58 == _GEN_9154 ? pht_7_88 : _GEN_1943; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1945 = 3'h7 == pht_rindex & 7'h59 == _GEN_9154 ? pht_7_89 : _GEN_1944; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1946 = 3'h7 == pht_rindex & 7'h5a == _GEN_9154 ? pht_7_90 : _GEN_1945; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1947 = 3'h7 == pht_rindex & 7'h5b == _GEN_9154 ? pht_7_91 : _GEN_1946; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1948 = 3'h7 == pht_rindex & 7'h5c == _GEN_9154 ? pht_7_92 : _GEN_1947; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1949 = 3'h7 == pht_rindex & 7'h5d == _GEN_9154 ? pht_7_93 : _GEN_1948; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1950 = 3'h7 == pht_rindex & 7'h5e == _GEN_9154 ? pht_7_94 : _GEN_1949; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1951 = 3'h7 == pht_rindex & 7'h5f == _GEN_9154 ? pht_7_95 : _GEN_1950; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1952 = 3'h7 == pht_rindex & 7'h60 == _GEN_9154 ? pht_7_96 : _GEN_1951; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1953 = 3'h7 == pht_rindex & 7'h61 == _GEN_9154 ? pht_7_97 : _GEN_1952; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1954 = 3'h7 == pht_rindex & 7'h62 == _GEN_9154 ? pht_7_98 : _GEN_1953; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1955 = 3'h7 == pht_rindex & 7'h63 == _GEN_9154 ? pht_7_99 : _GEN_1954; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1956 = 3'h7 == pht_rindex & 7'h64 == _GEN_9154 ? pht_7_100 : _GEN_1955; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1957 = 3'h7 == pht_rindex & 7'h65 == _GEN_9154 ? pht_7_101 : _GEN_1956; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1958 = 3'h7 == pht_rindex & 7'h66 == _GEN_9154 ? pht_7_102 : _GEN_1957; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1959 = 3'h7 == pht_rindex & 7'h67 == _GEN_9154 ? pht_7_103 : _GEN_1958; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1960 = 3'h7 == pht_rindex & 7'h68 == _GEN_9154 ? pht_7_104 : _GEN_1959; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1961 = 3'h7 == pht_rindex & 7'h69 == _GEN_9154 ? pht_7_105 : _GEN_1960; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1962 = 3'h7 == pht_rindex & 7'h6a == _GEN_9154 ? pht_7_106 : _GEN_1961; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1963 = 3'h7 == pht_rindex & 7'h6b == _GEN_9154 ? pht_7_107 : _GEN_1962; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1964 = 3'h7 == pht_rindex & 7'h6c == _GEN_9154 ? pht_7_108 : _GEN_1963; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1965 = 3'h7 == pht_rindex & 7'h6d == _GEN_9154 ? pht_7_109 : _GEN_1964; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1966 = 3'h7 == pht_rindex & 7'h6e == _GEN_9154 ? pht_7_110 : _GEN_1965; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1967 = 3'h7 == pht_rindex & 7'h6f == _GEN_9154 ? pht_7_111 : _GEN_1966; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1968 = 3'h7 == pht_rindex & 7'h70 == _GEN_9154 ? pht_7_112 : _GEN_1967; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1969 = 3'h7 == pht_rindex & 7'h71 == _GEN_9154 ? pht_7_113 : _GEN_1968; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1970 = 3'h7 == pht_rindex & 7'h72 == _GEN_9154 ? pht_7_114 : _GEN_1969; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1971 = 3'h7 == pht_rindex & 7'h73 == _GEN_9154 ? pht_7_115 : _GEN_1970; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1972 = 3'h7 == pht_rindex & 7'h74 == _GEN_9154 ? pht_7_116 : _GEN_1971; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1973 = 3'h7 == pht_rindex & 7'h75 == _GEN_9154 ? pht_7_117 : _GEN_1972; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1974 = 3'h7 == pht_rindex & 7'h76 == _GEN_9154 ? pht_7_118 : _GEN_1973; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1975 = 3'h7 == pht_rindex & 7'h77 == _GEN_9154 ? pht_7_119 : _GEN_1974; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1976 = 3'h7 == pht_rindex & 7'h78 == _GEN_9154 ? pht_7_120 : _GEN_1975; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1977 = 3'h7 == pht_rindex & 7'h79 == _GEN_9154 ? pht_7_121 : _GEN_1976; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1978 = 3'h7 == pht_rindex & 7'h7a == _GEN_9154 ? pht_7_122 : _GEN_1977; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1979 = 3'h7 == pht_rindex & 7'h7b == _GEN_9154 ? pht_7_123 : _GEN_1978; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1980 = 3'h7 == pht_rindex & 7'h7c == _GEN_9154 ? pht_7_124 : _GEN_1979; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1981 = 3'h7 == pht_rindex & 7'h7d == _GEN_9154 ? pht_7_125 : _GEN_1980; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1982 = 3'h7 == pht_rindex & 7'h7e == _GEN_9154 ? pht_7_126 : _GEN_1981; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1983 = 3'h7 == pht_rindex & 7'h7f == _GEN_9154 ? pht_7_127 : _GEN_1982; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1984 = 3'h7 == pht_rindex & 8'h80 == _GEN_9346 ? pht_7_128 : _GEN_1983; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1985 = 3'h7 == pht_rindex & 8'h81 == _GEN_9346 ? pht_7_129 : _GEN_1984; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1986 = 3'h7 == pht_rindex & 8'h82 == _GEN_9346 ? pht_7_130 : _GEN_1985; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1987 = 3'h7 == pht_rindex & 8'h83 == _GEN_9346 ? pht_7_131 : _GEN_1986; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1988 = 3'h7 == pht_rindex & 8'h84 == _GEN_9346 ? pht_7_132 : _GEN_1987; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1989 = 3'h7 == pht_rindex & 8'h85 == _GEN_9346 ? pht_7_133 : _GEN_1988; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1990 = 3'h7 == pht_rindex & 8'h86 == _GEN_9346 ? pht_7_134 : _GEN_1989; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1991 = 3'h7 == pht_rindex & 8'h87 == _GEN_9346 ? pht_7_135 : _GEN_1990; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1992 = 3'h7 == pht_rindex & 8'h88 == _GEN_9346 ? pht_7_136 : _GEN_1991; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1993 = 3'h7 == pht_rindex & 8'h89 == _GEN_9346 ? pht_7_137 : _GEN_1992; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1994 = 3'h7 == pht_rindex & 8'h8a == _GEN_9346 ? pht_7_138 : _GEN_1993; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1995 = 3'h7 == pht_rindex & 8'h8b == _GEN_9346 ? pht_7_139 : _GEN_1994; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1996 = 3'h7 == pht_rindex & 8'h8c == _GEN_9346 ? pht_7_140 : _GEN_1995; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1997 = 3'h7 == pht_rindex & 8'h8d == _GEN_9346 ? pht_7_141 : _GEN_1996; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1998 = 3'h7 == pht_rindex & 8'h8e == _GEN_9346 ? pht_7_142 : _GEN_1997; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_1999 = 3'h7 == pht_rindex & 8'h8f == _GEN_9346 ? pht_7_143 : _GEN_1998; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2000 = 3'h7 == pht_rindex & 8'h90 == _GEN_9346 ? pht_7_144 : _GEN_1999; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2001 = 3'h7 == pht_rindex & 8'h91 == _GEN_9346 ? pht_7_145 : _GEN_2000; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2002 = 3'h7 == pht_rindex & 8'h92 == _GEN_9346 ? pht_7_146 : _GEN_2001; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2003 = 3'h7 == pht_rindex & 8'h93 == _GEN_9346 ? pht_7_147 : _GEN_2002; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2004 = 3'h7 == pht_rindex & 8'h94 == _GEN_9346 ? pht_7_148 : _GEN_2003; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2005 = 3'h7 == pht_rindex & 8'h95 == _GEN_9346 ? pht_7_149 : _GEN_2004; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2006 = 3'h7 == pht_rindex & 8'h96 == _GEN_9346 ? pht_7_150 : _GEN_2005; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2007 = 3'h7 == pht_rindex & 8'h97 == _GEN_9346 ? pht_7_151 : _GEN_2006; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2008 = 3'h7 == pht_rindex & 8'h98 == _GEN_9346 ? pht_7_152 : _GEN_2007; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2009 = 3'h7 == pht_rindex & 8'h99 == _GEN_9346 ? pht_7_153 : _GEN_2008; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2010 = 3'h7 == pht_rindex & 8'h9a == _GEN_9346 ? pht_7_154 : _GEN_2009; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2011 = 3'h7 == pht_rindex & 8'h9b == _GEN_9346 ? pht_7_155 : _GEN_2010; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2012 = 3'h7 == pht_rindex & 8'h9c == _GEN_9346 ? pht_7_156 : _GEN_2011; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2013 = 3'h7 == pht_rindex & 8'h9d == _GEN_9346 ? pht_7_157 : _GEN_2012; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2014 = 3'h7 == pht_rindex & 8'h9e == _GEN_9346 ? pht_7_158 : _GEN_2013; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2015 = 3'h7 == pht_rindex & 8'h9f == _GEN_9346 ? pht_7_159 : _GEN_2014; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2016 = 3'h7 == pht_rindex & 8'ha0 == _GEN_9346 ? pht_7_160 : _GEN_2015; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2017 = 3'h7 == pht_rindex & 8'ha1 == _GEN_9346 ? pht_7_161 : _GEN_2016; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2018 = 3'h7 == pht_rindex & 8'ha2 == _GEN_9346 ? pht_7_162 : _GEN_2017; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2019 = 3'h7 == pht_rindex & 8'ha3 == _GEN_9346 ? pht_7_163 : _GEN_2018; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2020 = 3'h7 == pht_rindex & 8'ha4 == _GEN_9346 ? pht_7_164 : _GEN_2019; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2021 = 3'h7 == pht_rindex & 8'ha5 == _GEN_9346 ? pht_7_165 : _GEN_2020; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2022 = 3'h7 == pht_rindex & 8'ha6 == _GEN_9346 ? pht_7_166 : _GEN_2021; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2023 = 3'h7 == pht_rindex & 8'ha7 == _GEN_9346 ? pht_7_167 : _GEN_2022; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2024 = 3'h7 == pht_rindex & 8'ha8 == _GEN_9346 ? pht_7_168 : _GEN_2023; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2025 = 3'h7 == pht_rindex & 8'ha9 == _GEN_9346 ? pht_7_169 : _GEN_2024; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2026 = 3'h7 == pht_rindex & 8'haa == _GEN_9346 ? pht_7_170 : _GEN_2025; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2027 = 3'h7 == pht_rindex & 8'hab == _GEN_9346 ? pht_7_171 : _GEN_2026; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2028 = 3'h7 == pht_rindex & 8'hac == _GEN_9346 ? pht_7_172 : _GEN_2027; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2029 = 3'h7 == pht_rindex & 8'had == _GEN_9346 ? pht_7_173 : _GEN_2028; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2030 = 3'h7 == pht_rindex & 8'hae == _GEN_9346 ? pht_7_174 : _GEN_2029; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2031 = 3'h7 == pht_rindex & 8'haf == _GEN_9346 ? pht_7_175 : _GEN_2030; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2032 = 3'h7 == pht_rindex & 8'hb0 == _GEN_9346 ? pht_7_176 : _GEN_2031; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2033 = 3'h7 == pht_rindex & 8'hb1 == _GEN_9346 ? pht_7_177 : _GEN_2032; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2034 = 3'h7 == pht_rindex & 8'hb2 == _GEN_9346 ? pht_7_178 : _GEN_2033; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2035 = 3'h7 == pht_rindex & 8'hb3 == _GEN_9346 ? pht_7_179 : _GEN_2034; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2036 = 3'h7 == pht_rindex & 8'hb4 == _GEN_9346 ? pht_7_180 : _GEN_2035; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2037 = 3'h7 == pht_rindex & 8'hb5 == _GEN_9346 ? pht_7_181 : _GEN_2036; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2038 = 3'h7 == pht_rindex & 8'hb6 == _GEN_9346 ? pht_7_182 : _GEN_2037; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2039 = 3'h7 == pht_rindex & 8'hb7 == _GEN_9346 ? pht_7_183 : _GEN_2038; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2040 = 3'h7 == pht_rindex & 8'hb8 == _GEN_9346 ? pht_7_184 : _GEN_2039; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2041 = 3'h7 == pht_rindex & 8'hb9 == _GEN_9346 ? pht_7_185 : _GEN_2040; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2042 = 3'h7 == pht_rindex & 8'hba == _GEN_9346 ? pht_7_186 : _GEN_2041; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2043 = 3'h7 == pht_rindex & 8'hbb == _GEN_9346 ? pht_7_187 : _GEN_2042; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2044 = 3'h7 == pht_rindex & 8'hbc == _GEN_9346 ? pht_7_188 : _GEN_2043; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2045 = 3'h7 == pht_rindex & 8'hbd == _GEN_9346 ? pht_7_189 : _GEN_2044; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2046 = 3'h7 == pht_rindex & 8'hbe == _GEN_9346 ? pht_7_190 : _GEN_2045; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2047 = 3'h7 == pht_rindex & 8'hbf == _GEN_9346 ? pht_7_191 : _GEN_2046; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2048 = 3'h7 == pht_rindex & 8'hc0 == _GEN_9346 ? pht_7_192 : _GEN_2047; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2049 = 3'h7 == pht_rindex & 8'hc1 == _GEN_9346 ? pht_7_193 : _GEN_2048; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2050 = 3'h7 == pht_rindex & 8'hc2 == _GEN_9346 ? pht_7_194 : _GEN_2049; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2051 = 3'h7 == pht_rindex & 8'hc3 == _GEN_9346 ? pht_7_195 : _GEN_2050; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2052 = 3'h7 == pht_rindex & 8'hc4 == _GEN_9346 ? pht_7_196 : _GEN_2051; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2053 = 3'h7 == pht_rindex & 8'hc5 == _GEN_9346 ? pht_7_197 : _GEN_2052; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2054 = 3'h7 == pht_rindex & 8'hc6 == _GEN_9346 ? pht_7_198 : _GEN_2053; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2055 = 3'h7 == pht_rindex & 8'hc7 == _GEN_9346 ? pht_7_199 : _GEN_2054; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2056 = 3'h7 == pht_rindex & 8'hc8 == _GEN_9346 ? pht_7_200 : _GEN_2055; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2057 = 3'h7 == pht_rindex & 8'hc9 == _GEN_9346 ? pht_7_201 : _GEN_2056; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2058 = 3'h7 == pht_rindex & 8'hca == _GEN_9346 ? pht_7_202 : _GEN_2057; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2059 = 3'h7 == pht_rindex & 8'hcb == _GEN_9346 ? pht_7_203 : _GEN_2058; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2060 = 3'h7 == pht_rindex & 8'hcc == _GEN_9346 ? pht_7_204 : _GEN_2059; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2061 = 3'h7 == pht_rindex & 8'hcd == _GEN_9346 ? pht_7_205 : _GEN_2060; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2062 = 3'h7 == pht_rindex & 8'hce == _GEN_9346 ? pht_7_206 : _GEN_2061; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2063 = 3'h7 == pht_rindex & 8'hcf == _GEN_9346 ? pht_7_207 : _GEN_2062; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2064 = 3'h7 == pht_rindex & 8'hd0 == _GEN_9346 ? pht_7_208 : _GEN_2063; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2065 = 3'h7 == pht_rindex & 8'hd1 == _GEN_9346 ? pht_7_209 : _GEN_2064; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2066 = 3'h7 == pht_rindex & 8'hd2 == _GEN_9346 ? pht_7_210 : _GEN_2065; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2067 = 3'h7 == pht_rindex & 8'hd3 == _GEN_9346 ? pht_7_211 : _GEN_2066; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2068 = 3'h7 == pht_rindex & 8'hd4 == _GEN_9346 ? pht_7_212 : _GEN_2067; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2069 = 3'h7 == pht_rindex & 8'hd5 == _GEN_9346 ? pht_7_213 : _GEN_2068; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2070 = 3'h7 == pht_rindex & 8'hd6 == _GEN_9346 ? pht_7_214 : _GEN_2069; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2071 = 3'h7 == pht_rindex & 8'hd7 == _GEN_9346 ? pht_7_215 : _GEN_2070; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2072 = 3'h7 == pht_rindex & 8'hd8 == _GEN_9346 ? pht_7_216 : _GEN_2071; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2073 = 3'h7 == pht_rindex & 8'hd9 == _GEN_9346 ? pht_7_217 : _GEN_2072; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2074 = 3'h7 == pht_rindex & 8'hda == _GEN_9346 ? pht_7_218 : _GEN_2073; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2075 = 3'h7 == pht_rindex & 8'hdb == _GEN_9346 ? pht_7_219 : _GEN_2074; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2076 = 3'h7 == pht_rindex & 8'hdc == _GEN_9346 ? pht_7_220 : _GEN_2075; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2077 = 3'h7 == pht_rindex & 8'hdd == _GEN_9346 ? pht_7_221 : _GEN_2076; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2078 = 3'h7 == pht_rindex & 8'hde == _GEN_9346 ? pht_7_222 : _GEN_2077; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2079 = 3'h7 == pht_rindex & 8'hdf == _GEN_9346 ? pht_7_223 : _GEN_2078; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2080 = 3'h7 == pht_rindex & 8'he0 == _GEN_9346 ? pht_7_224 : _GEN_2079; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2081 = 3'h7 == pht_rindex & 8'he1 == _GEN_9346 ? pht_7_225 : _GEN_2080; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2082 = 3'h7 == pht_rindex & 8'he2 == _GEN_9346 ? pht_7_226 : _GEN_2081; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2083 = 3'h7 == pht_rindex & 8'he3 == _GEN_9346 ? pht_7_227 : _GEN_2082; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2084 = 3'h7 == pht_rindex & 8'he4 == _GEN_9346 ? pht_7_228 : _GEN_2083; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2085 = 3'h7 == pht_rindex & 8'he5 == _GEN_9346 ? pht_7_229 : _GEN_2084; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2086 = 3'h7 == pht_rindex & 8'he6 == _GEN_9346 ? pht_7_230 : _GEN_2085; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2087 = 3'h7 == pht_rindex & 8'he7 == _GEN_9346 ? pht_7_231 : _GEN_2086; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2088 = 3'h7 == pht_rindex & 8'he8 == _GEN_9346 ? pht_7_232 : _GEN_2087; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2089 = 3'h7 == pht_rindex & 8'he9 == _GEN_9346 ? pht_7_233 : _GEN_2088; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2090 = 3'h7 == pht_rindex & 8'hea == _GEN_9346 ? pht_7_234 : _GEN_2089; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2091 = 3'h7 == pht_rindex & 8'heb == _GEN_9346 ? pht_7_235 : _GEN_2090; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2092 = 3'h7 == pht_rindex & 8'hec == _GEN_9346 ? pht_7_236 : _GEN_2091; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2093 = 3'h7 == pht_rindex & 8'hed == _GEN_9346 ? pht_7_237 : _GEN_2092; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2094 = 3'h7 == pht_rindex & 8'hee == _GEN_9346 ? pht_7_238 : _GEN_2093; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2095 = 3'h7 == pht_rindex & 8'hef == _GEN_9346 ? pht_7_239 : _GEN_2094; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2096 = 3'h7 == pht_rindex & 8'hf0 == _GEN_9346 ? pht_7_240 : _GEN_2095; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2097 = 3'h7 == pht_rindex & 8'hf1 == _GEN_9346 ? pht_7_241 : _GEN_2096; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2098 = 3'h7 == pht_rindex & 8'hf2 == _GEN_9346 ? pht_7_242 : _GEN_2097; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2099 = 3'h7 == pht_rindex & 8'hf3 == _GEN_9346 ? pht_7_243 : _GEN_2098; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2100 = 3'h7 == pht_rindex & 8'hf4 == _GEN_9346 ? pht_7_244 : _GEN_2099; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2101 = 3'h7 == pht_rindex & 8'hf5 == _GEN_9346 ? pht_7_245 : _GEN_2100; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2102 = 3'h7 == pht_rindex & 8'hf6 == _GEN_9346 ? pht_7_246 : _GEN_2101; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2103 = 3'h7 == pht_rindex & 8'hf7 == _GEN_9346 ? pht_7_247 : _GEN_2102; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2104 = 3'h7 == pht_rindex & 8'hf8 == _GEN_9346 ? pht_7_248 : _GEN_2103; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2105 = 3'h7 == pht_rindex & 8'hf9 == _GEN_9346 ? pht_7_249 : _GEN_2104; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2106 = 3'h7 == pht_rindex & 8'hfa == _GEN_9346 ? pht_7_250 : _GEN_2105; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2107 = 3'h7 == pht_rindex & 8'hfb == _GEN_9346 ? pht_7_251 : _GEN_2106; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2108 = 3'h7 == pht_rindex & 8'hfc == _GEN_9346 ? pht_7_252 : _GEN_2107; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2109 = 3'h7 == pht_rindex & 8'hfd == _GEN_9346 ? pht_7_253 : _GEN_2108; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2110 = 3'h7 == pht_rindex & 8'hfe == _GEN_9346 ? pht_7_254 : _GEN_2109; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire [1:0] _GEN_2111 = 3'h7 == pht_rindex & 8'hff == _GEN_9346 ? pht_7_255 : _GEN_2110; // @[BrPredictor.scala 62:47 BrPredictor.scala 62:47]
  wire  pht_rdirect = _GEN_2111[1]; // @[BrPredictor.scala 62:47]
  wire [5:0] bht_waddr = io_jmp_packet_inst_pc[7:2]; // @[BrPredictor.scala 52:34]
  wire [5:0] _GEN_2113 = 6'h1 == bht_waddr ? bht_1 : bht_0; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2114 = 6'h2 == bht_waddr ? bht_2 : _GEN_2113; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2115 = 6'h3 == bht_waddr ? bht_3 : _GEN_2114; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2116 = 6'h4 == bht_waddr ? bht_4 : _GEN_2115; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2117 = 6'h5 == bht_waddr ? bht_5 : _GEN_2116; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2118 = 6'h6 == bht_waddr ? bht_6 : _GEN_2117; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2119 = 6'h7 == bht_waddr ? bht_7 : _GEN_2118; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2120 = 6'h8 == bht_waddr ? bht_8 : _GEN_2119; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2121 = 6'h9 == bht_waddr ? bht_9 : _GEN_2120; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2122 = 6'ha == bht_waddr ? bht_10 : _GEN_2121; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2123 = 6'hb == bht_waddr ? bht_11 : _GEN_2122; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2124 = 6'hc == bht_waddr ? bht_12 : _GEN_2123; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2125 = 6'hd == bht_waddr ? bht_13 : _GEN_2124; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2126 = 6'he == bht_waddr ? bht_14 : _GEN_2125; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2127 = 6'hf == bht_waddr ? bht_15 : _GEN_2126; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2128 = 6'h10 == bht_waddr ? bht_16 : _GEN_2127; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2129 = 6'h11 == bht_waddr ? bht_17 : _GEN_2128; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2130 = 6'h12 == bht_waddr ? bht_18 : _GEN_2129; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2131 = 6'h13 == bht_waddr ? bht_19 : _GEN_2130; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2132 = 6'h14 == bht_waddr ? bht_20 : _GEN_2131; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2133 = 6'h15 == bht_waddr ? bht_21 : _GEN_2132; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2134 = 6'h16 == bht_waddr ? bht_22 : _GEN_2133; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2135 = 6'h17 == bht_waddr ? bht_23 : _GEN_2134; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2136 = 6'h18 == bht_waddr ? bht_24 : _GEN_2135; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2137 = 6'h19 == bht_waddr ? bht_25 : _GEN_2136; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2138 = 6'h1a == bht_waddr ? bht_26 : _GEN_2137; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2139 = 6'h1b == bht_waddr ? bht_27 : _GEN_2138; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2140 = 6'h1c == bht_waddr ? bht_28 : _GEN_2139; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2141 = 6'h1d == bht_waddr ? bht_29 : _GEN_2140; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2142 = 6'h1e == bht_waddr ? bht_30 : _GEN_2141; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2143 = 6'h1f == bht_waddr ? bht_31 : _GEN_2142; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2144 = 6'h20 == bht_waddr ? bht_32 : _GEN_2143; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2145 = 6'h21 == bht_waddr ? bht_33 : _GEN_2144; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2146 = 6'h22 == bht_waddr ? bht_34 : _GEN_2145; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2147 = 6'h23 == bht_waddr ? bht_35 : _GEN_2146; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2148 = 6'h24 == bht_waddr ? bht_36 : _GEN_2147; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2149 = 6'h25 == bht_waddr ? bht_37 : _GEN_2148; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2150 = 6'h26 == bht_waddr ? bht_38 : _GEN_2149; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2151 = 6'h27 == bht_waddr ? bht_39 : _GEN_2150; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2152 = 6'h28 == bht_waddr ? bht_40 : _GEN_2151; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2153 = 6'h29 == bht_waddr ? bht_41 : _GEN_2152; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2154 = 6'h2a == bht_waddr ? bht_42 : _GEN_2153; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2155 = 6'h2b == bht_waddr ? bht_43 : _GEN_2154; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2156 = 6'h2c == bht_waddr ? bht_44 : _GEN_2155; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2157 = 6'h2d == bht_waddr ? bht_45 : _GEN_2156; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2158 = 6'h2e == bht_waddr ? bht_46 : _GEN_2157; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2159 = 6'h2f == bht_waddr ? bht_47 : _GEN_2158; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2160 = 6'h30 == bht_waddr ? bht_48 : _GEN_2159; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2161 = 6'h31 == bht_waddr ? bht_49 : _GEN_2160; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2162 = 6'h32 == bht_waddr ? bht_50 : _GEN_2161; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2163 = 6'h33 == bht_waddr ? bht_51 : _GEN_2162; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2164 = 6'h34 == bht_waddr ? bht_52 : _GEN_2163; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2165 = 6'h35 == bht_waddr ? bht_53 : _GEN_2164; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2166 = 6'h36 == bht_waddr ? bht_54 : _GEN_2165; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2167 = 6'h37 == bht_waddr ? bht_55 : _GEN_2166; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2168 = 6'h38 == bht_waddr ? bht_56 : _GEN_2167; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2169 = 6'h39 == bht_waddr ? bht_57 : _GEN_2168; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2170 = 6'h3a == bht_waddr ? bht_58 : _GEN_2169; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2171 = 6'h3b == bht_waddr ? bht_59 : _GEN_2170; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2172 = 6'h3c == bht_waddr ? bht_60 : _GEN_2171; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2173 = 6'h3d == bht_waddr ? bht_61 : _GEN_2172; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2174 = 6'h3e == bht_waddr ? bht_62 : _GEN_2173; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [5:0] _GEN_2175 = 6'h3f == bht_waddr ? bht_63 : _GEN_2174; // @[BrPredictor.scala 69:62 BrPredictor.scala 69:62]
  wire [4:0] bht_lo = _GEN_2175[5:1]; // @[BrPredictor.scala 69:62]
  wire [5:0] _bht_T = {io_jmp_packet_jmp,bht_lo}; // @[Cat.scala 30:58]
  wire [5:0] pht_waddr = _GEN_2175 ^ bht_waddr; // @[BrPredictor.scala 53:58]
  wire [2:0] pht_windex = io_jmp_packet_inst_pc[10:8]; // @[BrPredictor.scala 54:35]
  wire [1:0] _pht_T_1 = io_jmp_packet_jmp ? 2'h2 : 2'h0; // @[BrPredictor.scala 77:17]
  wire [1:0] _pht_T_2 = io_jmp_packet_jmp ? 2'h3 : 2'h1; // @[BrPredictor.scala 78:17]
  wire [1:0] _pht_T_3 = io_jmp_packet_jmp ? 2'h3 : 2'h2; // @[BrPredictor.scala 79:17]
  wire  _GEN_14658 = 3'h0 == pht_windex; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14659 = 6'h1 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2305 = 3'h0 == pht_windex & 6'h1 == pht_waddr ? pht_0_1 : pht_0_0; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14661 = 6'h2 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2306 = 3'h0 == pht_windex & 6'h2 == pht_waddr ? pht_0_2 : _GEN_2305; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14663 = 6'h3 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2307 = 3'h0 == pht_windex & 6'h3 == pht_waddr ? pht_0_3 : _GEN_2306; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14665 = 6'h4 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2308 = 3'h0 == pht_windex & 6'h4 == pht_waddr ? pht_0_4 : _GEN_2307; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14667 = 6'h5 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2309 = 3'h0 == pht_windex & 6'h5 == pht_waddr ? pht_0_5 : _GEN_2308; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14669 = 6'h6 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2310 = 3'h0 == pht_windex & 6'h6 == pht_waddr ? pht_0_6 : _GEN_2309; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14671 = 6'h7 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2311 = 3'h0 == pht_windex & 6'h7 == pht_waddr ? pht_0_7 : _GEN_2310; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14673 = 6'h8 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2312 = 3'h0 == pht_windex & 6'h8 == pht_waddr ? pht_0_8 : _GEN_2311; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14675 = 6'h9 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2313 = 3'h0 == pht_windex & 6'h9 == pht_waddr ? pht_0_9 : _GEN_2312; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14677 = 6'ha == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2314 = 3'h0 == pht_windex & 6'ha == pht_waddr ? pht_0_10 : _GEN_2313; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14679 = 6'hb == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2315 = 3'h0 == pht_windex & 6'hb == pht_waddr ? pht_0_11 : _GEN_2314; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14681 = 6'hc == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2316 = 3'h0 == pht_windex & 6'hc == pht_waddr ? pht_0_12 : _GEN_2315; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14683 = 6'hd == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2317 = 3'h0 == pht_windex & 6'hd == pht_waddr ? pht_0_13 : _GEN_2316; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14685 = 6'he == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2318 = 3'h0 == pht_windex & 6'he == pht_waddr ? pht_0_14 : _GEN_2317; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14687 = 6'hf == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2319 = 3'h0 == pht_windex & 6'hf == pht_waddr ? pht_0_15 : _GEN_2318; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14689 = 6'h10 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2320 = 3'h0 == pht_windex & 6'h10 == pht_waddr ? pht_0_16 : _GEN_2319; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14691 = 6'h11 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2321 = 3'h0 == pht_windex & 6'h11 == pht_waddr ? pht_0_17 : _GEN_2320; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14693 = 6'h12 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2322 = 3'h0 == pht_windex & 6'h12 == pht_waddr ? pht_0_18 : _GEN_2321; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14695 = 6'h13 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2323 = 3'h0 == pht_windex & 6'h13 == pht_waddr ? pht_0_19 : _GEN_2322; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14697 = 6'h14 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2324 = 3'h0 == pht_windex & 6'h14 == pht_waddr ? pht_0_20 : _GEN_2323; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14699 = 6'h15 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2325 = 3'h0 == pht_windex & 6'h15 == pht_waddr ? pht_0_21 : _GEN_2324; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14701 = 6'h16 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2326 = 3'h0 == pht_windex & 6'h16 == pht_waddr ? pht_0_22 : _GEN_2325; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14703 = 6'h17 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2327 = 3'h0 == pht_windex & 6'h17 == pht_waddr ? pht_0_23 : _GEN_2326; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14705 = 6'h18 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2328 = 3'h0 == pht_windex & 6'h18 == pht_waddr ? pht_0_24 : _GEN_2327; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14707 = 6'h19 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2329 = 3'h0 == pht_windex & 6'h19 == pht_waddr ? pht_0_25 : _GEN_2328; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14709 = 6'h1a == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2330 = 3'h0 == pht_windex & 6'h1a == pht_waddr ? pht_0_26 : _GEN_2329; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14711 = 6'h1b == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2331 = 3'h0 == pht_windex & 6'h1b == pht_waddr ? pht_0_27 : _GEN_2330; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14713 = 6'h1c == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2332 = 3'h0 == pht_windex & 6'h1c == pht_waddr ? pht_0_28 : _GEN_2331; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14715 = 6'h1d == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2333 = 3'h0 == pht_windex & 6'h1d == pht_waddr ? pht_0_29 : _GEN_2332; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14717 = 6'h1e == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2334 = 3'h0 == pht_windex & 6'h1e == pht_waddr ? pht_0_30 : _GEN_2333; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14719 = 6'h1f == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2335 = 3'h0 == pht_windex & 6'h1f == pht_waddr ? pht_0_31 : _GEN_2334; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14721 = 6'h20 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2336 = 3'h0 == pht_windex & 6'h20 == pht_waddr ? pht_0_32 : _GEN_2335; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14723 = 6'h21 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2337 = 3'h0 == pht_windex & 6'h21 == pht_waddr ? pht_0_33 : _GEN_2336; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14725 = 6'h22 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2338 = 3'h0 == pht_windex & 6'h22 == pht_waddr ? pht_0_34 : _GEN_2337; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14727 = 6'h23 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2339 = 3'h0 == pht_windex & 6'h23 == pht_waddr ? pht_0_35 : _GEN_2338; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14729 = 6'h24 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2340 = 3'h0 == pht_windex & 6'h24 == pht_waddr ? pht_0_36 : _GEN_2339; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14731 = 6'h25 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2341 = 3'h0 == pht_windex & 6'h25 == pht_waddr ? pht_0_37 : _GEN_2340; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14733 = 6'h26 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2342 = 3'h0 == pht_windex & 6'h26 == pht_waddr ? pht_0_38 : _GEN_2341; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14735 = 6'h27 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2343 = 3'h0 == pht_windex & 6'h27 == pht_waddr ? pht_0_39 : _GEN_2342; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14737 = 6'h28 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2344 = 3'h0 == pht_windex & 6'h28 == pht_waddr ? pht_0_40 : _GEN_2343; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14739 = 6'h29 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2345 = 3'h0 == pht_windex & 6'h29 == pht_waddr ? pht_0_41 : _GEN_2344; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14741 = 6'h2a == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2346 = 3'h0 == pht_windex & 6'h2a == pht_waddr ? pht_0_42 : _GEN_2345; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14743 = 6'h2b == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2347 = 3'h0 == pht_windex & 6'h2b == pht_waddr ? pht_0_43 : _GEN_2346; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14745 = 6'h2c == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2348 = 3'h0 == pht_windex & 6'h2c == pht_waddr ? pht_0_44 : _GEN_2347; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14747 = 6'h2d == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2349 = 3'h0 == pht_windex & 6'h2d == pht_waddr ? pht_0_45 : _GEN_2348; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14749 = 6'h2e == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2350 = 3'h0 == pht_windex & 6'h2e == pht_waddr ? pht_0_46 : _GEN_2349; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14751 = 6'h2f == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2351 = 3'h0 == pht_windex & 6'h2f == pht_waddr ? pht_0_47 : _GEN_2350; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14753 = 6'h30 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2352 = 3'h0 == pht_windex & 6'h30 == pht_waddr ? pht_0_48 : _GEN_2351; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14755 = 6'h31 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2353 = 3'h0 == pht_windex & 6'h31 == pht_waddr ? pht_0_49 : _GEN_2352; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14757 = 6'h32 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2354 = 3'h0 == pht_windex & 6'h32 == pht_waddr ? pht_0_50 : _GEN_2353; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14759 = 6'h33 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2355 = 3'h0 == pht_windex & 6'h33 == pht_waddr ? pht_0_51 : _GEN_2354; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14761 = 6'h34 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2356 = 3'h0 == pht_windex & 6'h34 == pht_waddr ? pht_0_52 : _GEN_2355; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14763 = 6'h35 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2357 = 3'h0 == pht_windex & 6'h35 == pht_waddr ? pht_0_53 : _GEN_2356; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14765 = 6'h36 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2358 = 3'h0 == pht_windex & 6'h36 == pht_waddr ? pht_0_54 : _GEN_2357; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14767 = 6'h37 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2359 = 3'h0 == pht_windex & 6'h37 == pht_waddr ? pht_0_55 : _GEN_2358; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14769 = 6'h38 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2360 = 3'h0 == pht_windex & 6'h38 == pht_waddr ? pht_0_56 : _GEN_2359; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14771 = 6'h39 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2361 = 3'h0 == pht_windex & 6'h39 == pht_waddr ? pht_0_57 : _GEN_2360; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14773 = 6'h3a == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2362 = 3'h0 == pht_windex & 6'h3a == pht_waddr ? pht_0_58 : _GEN_2361; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14775 = 6'h3b == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2363 = 3'h0 == pht_windex & 6'h3b == pht_waddr ? pht_0_59 : _GEN_2362; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14777 = 6'h3c == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2364 = 3'h0 == pht_windex & 6'h3c == pht_waddr ? pht_0_60 : _GEN_2363; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14779 = 6'h3d == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2365 = 3'h0 == pht_windex & 6'h3d == pht_waddr ? pht_0_61 : _GEN_2364; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14781 = 6'h3e == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2366 = 3'h0 == pht_windex & 6'h3e == pht_waddr ? pht_0_62 : _GEN_2365; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14783 = 6'h3f == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2367 = 3'h0 == pht_windex & 6'h3f == pht_waddr ? pht_0_63 : _GEN_2366; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [6:0] _GEN_14784 = {{1'd0}, pht_waddr}; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14786 = 7'h40 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2368 = 3'h0 == pht_windex & 7'h40 == _GEN_14784 ? pht_0_64 : _GEN_2367; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14789 = 7'h41 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2369 = 3'h0 == pht_windex & 7'h41 == _GEN_14784 ? pht_0_65 : _GEN_2368; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14792 = 7'h42 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2370 = 3'h0 == pht_windex & 7'h42 == _GEN_14784 ? pht_0_66 : _GEN_2369; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14795 = 7'h43 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2371 = 3'h0 == pht_windex & 7'h43 == _GEN_14784 ? pht_0_67 : _GEN_2370; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14798 = 7'h44 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2372 = 3'h0 == pht_windex & 7'h44 == _GEN_14784 ? pht_0_68 : _GEN_2371; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14801 = 7'h45 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2373 = 3'h0 == pht_windex & 7'h45 == _GEN_14784 ? pht_0_69 : _GEN_2372; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14804 = 7'h46 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2374 = 3'h0 == pht_windex & 7'h46 == _GEN_14784 ? pht_0_70 : _GEN_2373; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14807 = 7'h47 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2375 = 3'h0 == pht_windex & 7'h47 == _GEN_14784 ? pht_0_71 : _GEN_2374; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14810 = 7'h48 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2376 = 3'h0 == pht_windex & 7'h48 == _GEN_14784 ? pht_0_72 : _GEN_2375; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14813 = 7'h49 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2377 = 3'h0 == pht_windex & 7'h49 == _GEN_14784 ? pht_0_73 : _GEN_2376; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14816 = 7'h4a == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2378 = 3'h0 == pht_windex & 7'h4a == _GEN_14784 ? pht_0_74 : _GEN_2377; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14819 = 7'h4b == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2379 = 3'h0 == pht_windex & 7'h4b == _GEN_14784 ? pht_0_75 : _GEN_2378; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14822 = 7'h4c == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2380 = 3'h0 == pht_windex & 7'h4c == _GEN_14784 ? pht_0_76 : _GEN_2379; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14825 = 7'h4d == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2381 = 3'h0 == pht_windex & 7'h4d == _GEN_14784 ? pht_0_77 : _GEN_2380; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14828 = 7'h4e == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2382 = 3'h0 == pht_windex & 7'h4e == _GEN_14784 ? pht_0_78 : _GEN_2381; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14831 = 7'h4f == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2383 = 3'h0 == pht_windex & 7'h4f == _GEN_14784 ? pht_0_79 : _GEN_2382; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14834 = 7'h50 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2384 = 3'h0 == pht_windex & 7'h50 == _GEN_14784 ? pht_0_80 : _GEN_2383; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14837 = 7'h51 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2385 = 3'h0 == pht_windex & 7'h51 == _GEN_14784 ? pht_0_81 : _GEN_2384; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14840 = 7'h52 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2386 = 3'h0 == pht_windex & 7'h52 == _GEN_14784 ? pht_0_82 : _GEN_2385; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14843 = 7'h53 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2387 = 3'h0 == pht_windex & 7'h53 == _GEN_14784 ? pht_0_83 : _GEN_2386; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14846 = 7'h54 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2388 = 3'h0 == pht_windex & 7'h54 == _GEN_14784 ? pht_0_84 : _GEN_2387; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14849 = 7'h55 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2389 = 3'h0 == pht_windex & 7'h55 == _GEN_14784 ? pht_0_85 : _GEN_2388; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14852 = 7'h56 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2390 = 3'h0 == pht_windex & 7'h56 == _GEN_14784 ? pht_0_86 : _GEN_2389; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14855 = 7'h57 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2391 = 3'h0 == pht_windex & 7'h57 == _GEN_14784 ? pht_0_87 : _GEN_2390; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14858 = 7'h58 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2392 = 3'h0 == pht_windex & 7'h58 == _GEN_14784 ? pht_0_88 : _GEN_2391; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14861 = 7'h59 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2393 = 3'h0 == pht_windex & 7'h59 == _GEN_14784 ? pht_0_89 : _GEN_2392; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14864 = 7'h5a == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2394 = 3'h0 == pht_windex & 7'h5a == _GEN_14784 ? pht_0_90 : _GEN_2393; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14867 = 7'h5b == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2395 = 3'h0 == pht_windex & 7'h5b == _GEN_14784 ? pht_0_91 : _GEN_2394; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14870 = 7'h5c == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2396 = 3'h0 == pht_windex & 7'h5c == _GEN_14784 ? pht_0_92 : _GEN_2395; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14873 = 7'h5d == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2397 = 3'h0 == pht_windex & 7'h5d == _GEN_14784 ? pht_0_93 : _GEN_2396; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14876 = 7'h5e == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2398 = 3'h0 == pht_windex & 7'h5e == _GEN_14784 ? pht_0_94 : _GEN_2397; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14879 = 7'h5f == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2399 = 3'h0 == pht_windex & 7'h5f == _GEN_14784 ? pht_0_95 : _GEN_2398; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14882 = 7'h60 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2400 = 3'h0 == pht_windex & 7'h60 == _GEN_14784 ? pht_0_96 : _GEN_2399; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14885 = 7'h61 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2401 = 3'h0 == pht_windex & 7'h61 == _GEN_14784 ? pht_0_97 : _GEN_2400; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14888 = 7'h62 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2402 = 3'h0 == pht_windex & 7'h62 == _GEN_14784 ? pht_0_98 : _GEN_2401; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14891 = 7'h63 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2403 = 3'h0 == pht_windex & 7'h63 == _GEN_14784 ? pht_0_99 : _GEN_2402; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14894 = 7'h64 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2404 = 3'h0 == pht_windex & 7'h64 == _GEN_14784 ? pht_0_100 : _GEN_2403; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14897 = 7'h65 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2405 = 3'h0 == pht_windex & 7'h65 == _GEN_14784 ? pht_0_101 : _GEN_2404; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14900 = 7'h66 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2406 = 3'h0 == pht_windex & 7'h66 == _GEN_14784 ? pht_0_102 : _GEN_2405; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14903 = 7'h67 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2407 = 3'h0 == pht_windex & 7'h67 == _GEN_14784 ? pht_0_103 : _GEN_2406; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14906 = 7'h68 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2408 = 3'h0 == pht_windex & 7'h68 == _GEN_14784 ? pht_0_104 : _GEN_2407; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14909 = 7'h69 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2409 = 3'h0 == pht_windex & 7'h69 == _GEN_14784 ? pht_0_105 : _GEN_2408; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14912 = 7'h6a == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2410 = 3'h0 == pht_windex & 7'h6a == _GEN_14784 ? pht_0_106 : _GEN_2409; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14915 = 7'h6b == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2411 = 3'h0 == pht_windex & 7'h6b == _GEN_14784 ? pht_0_107 : _GEN_2410; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14918 = 7'h6c == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2412 = 3'h0 == pht_windex & 7'h6c == _GEN_14784 ? pht_0_108 : _GEN_2411; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14921 = 7'h6d == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2413 = 3'h0 == pht_windex & 7'h6d == _GEN_14784 ? pht_0_109 : _GEN_2412; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14924 = 7'h6e == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2414 = 3'h0 == pht_windex & 7'h6e == _GEN_14784 ? pht_0_110 : _GEN_2413; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14927 = 7'h6f == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2415 = 3'h0 == pht_windex & 7'h6f == _GEN_14784 ? pht_0_111 : _GEN_2414; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14930 = 7'h70 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2416 = 3'h0 == pht_windex & 7'h70 == _GEN_14784 ? pht_0_112 : _GEN_2415; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14933 = 7'h71 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2417 = 3'h0 == pht_windex & 7'h71 == _GEN_14784 ? pht_0_113 : _GEN_2416; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14936 = 7'h72 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2418 = 3'h0 == pht_windex & 7'h72 == _GEN_14784 ? pht_0_114 : _GEN_2417; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14939 = 7'h73 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2419 = 3'h0 == pht_windex & 7'h73 == _GEN_14784 ? pht_0_115 : _GEN_2418; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14942 = 7'h74 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2420 = 3'h0 == pht_windex & 7'h74 == _GEN_14784 ? pht_0_116 : _GEN_2419; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14945 = 7'h75 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2421 = 3'h0 == pht_windex & 7'h75 == _GEN_14784 ? pht_0_117 : _GEN_2420; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14948 = 7'h76 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2422 = 3'h0 == pht_windex & 7'h76 == _GEN_14784 ? pht_0_118 : _GEN_2421; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14951 = 7'h77 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2423 = 3'h0 == pht_windex & 7'h77 == _GEN_14784 ? pht_0_119 : _GEN_2422; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14954 = 7'h78 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2424 = 3'h0 == pht_windex & 7'h78 == _GEN_14784 ? pht_0_120 : _GEN_2423; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14957 = 7'h79 == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2425 = 3'h0 == pht_windex & 7'h79 == _GEN_14784 ? pht_0_121 : _GEN_2424; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14960 = 7'h7a == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2426 = 3'h0 == pht_windex & 7'h7a == _GEN_14784 ? pht_0_122 : _GEN_2425; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14963 = 7'h7b == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2427 = 3'h0 == pht_windex & 7'h7b == _GEN_14784 ? pht_0_123 : _GEN_2426; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14966 = 7'h7c == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2428 = 3'h0 == pht_windex & 7'h7c == _GEN_14784 ? pht_0_124 : _GEN_2427; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14969 = 7'h7d == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2429 = 3'h0 == pht_windex & 7'h7d == _GEN_14784 ? pht_0_125 : _GEN_2428; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14972 = 7'h7e == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2430 = 3'h0 == pht_windex & 7'h7e == _GEN_14784 ? pht_0_126 : _GEN_2429; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14975 = 7'h7f == _GEN_14784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2431 = 3'h0 == pht_windex & 7'h7f == _GEN_14784 ? pht_0_127 : _GEN_2430; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [7:0] _GEN_14976 = {{2'd0}, pht_waddr}; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14978 = 8'h80 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2432 = 3'h0 == pht_windex & 8'h80 == _GEN_14976 ? pht_0_128 : _GEN_2431; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14981 = 8'h81 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2433 = 3'h0 == pht_windex & 8'h81 == _GEN_14976 ? pht_0_129 : _GEN_2432; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14984 = 8'h82 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2434 = 3'h0 == pht_windex & 8'h82 == _GEN_14976 ? pht_0_130 : _GEN_2433; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14987 = 8'h83 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2435 = 3'h0 == pht_windex & 8'h83 == _GEN_14976 ? pht_0_131 : _GEN_2434; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14990 = 8'h84 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2436 = 3'h0 == pht_windex & 8'h84 == _GEN_14976 ? pht_0_132 : _GEN_2435; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14993 = 8'h85 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2437 = 3'h0 == pht_windex & 8'h85 == _GEN_14976 ? pht_0_133 : _GEN_2436; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14996 = 8'h86 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2438 = 3'h0 == pht_windex & 8'h86 == _GEN_14976 ? pht_0_134 : _GEN_2437; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_14999 = 8'h87 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2439 = 3'h0 == pht_windex & 8'h87 == _GEN_14976 ? pht_0_135 : _GEN_2438; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15002 = 8'h88 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2440 = 3'h0 == pht_windex & 8'h88 == _GEN_14976 ? pht_0_136 : _GEN_2439; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15005 = 8'h89 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2441 = 3'h0 == pht_windex & 8'h89 == _GEN_14976 ? pht_0_137 : _GEN_2440; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15008 = 8'h8a == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2442 = 3'h0 == pht_windex & 8'h8a == _GEN_14976 ? pht_0_138 : _GEN_2441; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15011 = 8'h8b == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2443 = 3'h0 == pht_windex & 8'h8b == _GEN_14976 ? pht_0_139 : _GEN_2442; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15014 = 8'h8c == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2444 = 3'h0 == pht_windex & 8'h8c == _GEN_14976 ? pht_0_140 : _GEN_2443; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15017 = 8'h8d == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2445 = 3'h0 == pht_windex & 8'h8d == _GEN_14976 ? pht_0_141 : _GEN_2444; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15020 = 8'h8e == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2446 = 3'h0 == pht_windex & 8'h8e == _GEN_14976 ? pht_0_142 : _GEN_2445; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15023 = 8'h8f == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2447 = 3'h0 == pht_windex & 8'h8f == _GEN_14976 ? pht_0_143 : _GEN_2446; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15026 = 8'h90 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2448 = 3'h0 == pht_windex & 8'h90 == _GEN_14976 ? pht_0_144 : _GEN_2447; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15029 = 8'h91 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2449 = 3'h0 == pht_windex & 8'h91 == _GEN_14976 ? pht_0_145 : _GEN_2448; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15032 = 8'h92 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2450 = 3'h0 == pht_windex & 8'h92 == _GEN_14976 ? pht_0_146 : _GEN_2449; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15035 = 8'h93 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2451 = 3'h0 == pht_windex & 8'h93 == _GEN_14976 ? pht_0_147 : _GEN_2450; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15038 = 8'h94 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2452 = 3'h0 == pht_windex & 8'h94 == _GEN_14976 ? pht_0_148 : _GEN_2451; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15041 = 8'h95 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2453 = 3'h0 == pht_windex & 8'h95 == _GEN_14976 ? pht_0_149 : _GEN_2452; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15044 = 8'h96 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2454 = 3'h0 == pht_windex & 8'h96 == _GEN_14976 ? pht_0_150 : _GEN_2453; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15047 = 8'h97 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2455 = 3'h0 == pht_windex & 8'h97 == _GEN_14976 ? pht_0_151 : _GEN_2454; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15050 = 8'h98 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2456 = 3'h0 == pht_windex & 8'h98 == _GEN_14976 ? pht_0_152 : _GEN_2455; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15053 = 8'h99 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2457 = 3'h0 == pht_windex & 8'h99 == _GEN_14976 ? pht_0_153 : _GEN_2456; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15056 = 8'h9a == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2458 = 3'h0 == pht_windex & 8'h9a == _GEN_14976 ? pht_0_154 : _GEN_2457; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15059 = 8'h9b == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2459 = 3'h0 == pht_windex & 8'h9b == _GEN_14976 ? pht_0_155 : _GEN_2458; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15062 = 8'h9c == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2460 = 3'h0 == pht_windex & 8'h9c == _GEN_14976 ? pht_0_156 : _GEN_2459; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15065 = 8'h9d == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2461 = 3'h0 == pht_windex & 8'h9d == _GEN_14976 ? pht_0_157 : _GEN_2460; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15068 = 8'h9e == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2462 = 3'h0 == pht_windex & 8'h9e == _GEN_14976 ? pht_0_158 : _GEN_2461; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15071 = 8'h9f == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2463 = 3'h0 == pht_windex & 8'h9f == _GEN_14976 ? pht_0_159 : _GEN_2462; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15074 = 8'ha0 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2464 = 3'h0 == pht_windex & 8'ha0 == _GEN_14976 ? pht_0_160 : _GEN_2463; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15077 = 8'ha1 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2465 = 3'h0 == pht_windex & 8'ha1 == _GEN_14976 ? pht_0_161 : _GEN_2464; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15080 = 8'ha2 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2466 = 3'h0 == pht_windex & 8'ha2 == _GEN_14976 ? pht_0_162 : _GEN_2465; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15083 = 8'ha3 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2467 = 3'h0 == pht_windex & 8'ha3 == _GEN_14976 ? pht_0_163 : _GEN_2466; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15086 = 8'ha4 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2468 = 3'h0 == pht_windex & 8'ha4 == _GEN_14976 ? pht_0_164 : _GEN_2467; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15089 = 8'ha5 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2469 = 3'h0 == pht_windex & 8'ha5 == _GEN_14976 ? pht_0_165 : _GEN_2468; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15092 = 8'ha6 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2470 = 3'h0 == pht_windex & 8'ha6 == _GEN_14976 ? pht_0_166 : _GEN_2469; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15095 = 8'ha7 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2471 = 3'h0 == pht_windex & 8'ha7 == _GEN_14976 ? pht_0_167 : _GEN_2470; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15098 = 8'ha8 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2472 = 3'h0 == pht_windex & 8'ha8 == _GEN_14976 ? pht_0_168 : _GEN_2471; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15101 = 8'ha9 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2473 = 3'h0 == pht_windex & 8'ha9 == _GEN_14976 ? pht_0_169 : _GEN_2472; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15104 = 8'haa == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2474 = 3'h0 == pht_windex & 8'haa == _GEN_14976 ? pht_0_170 : _GEN_2473; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15107 = 8'hab == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2475 = 3'h0 == pht_windex & 8'hab == _GEN_14976 ? pht_0_171 : _GEN_2474; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15110 = 8'hac == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2476 = 3'h0 == pht_windex & 8'hac == _GEN_14976 ? pht_0_172 : _GEN_2475; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15113 = 8'had == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2477 = 3'h0 == pht_windex & 8'had == _GEN_14976 ? pht_0_173 : _GEN_2476; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15116 = 8'hae == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2478 = 3'h0 == pht_windex & 8'hae == _GEN_14976 ? pht_0_174 : _GEN_2477; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15119 = 8'haf == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2479 = 3'h0 == pht_windex & 8'haf == _GEN_14976 ? pht_0_175 : _GEN_2478; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15122 = 8'hb0 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2480 = 3'h0 == pht_windex & 8'hb0 == _GEN_14976 ? pht_0_176 : _GEN_2479; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15125 = 8'hb1 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2481 = 3'h0 == pht_windex & 8'hb1 == _GEN_14976 ? pht_0_177 : _GEN_2480; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15128 = 8'hb2 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2482 = 3'h0 == pht_windex & 8'hb2 == _GEN_14976 ? pht_0_178 : _GEN_2481; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15131 = 8'hb3 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2483 = 3'h0 == pht_windex & 8'hb3 == _GEN_14976 ? pht_0_179 : _GEN_2482; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15134 = 8'hb4 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2484 = 3'h0 == pht_windex & 8'hb4 == _GEN_14976 ? pht_0_180 : _GEN_2483; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15137 = 8'hb5 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2485 = 3'h0 == pht_windex & 8'hb5 == _GEN_14976 ? pht_0_181 : _GEN_2484; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15140 = 8'hb6 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2486 = 3'h0 == pht_windex & 8'hb6 == _GEN_14976 ? pht_0_182 : _GEN_2485; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15143 = 8'hb7 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2487 = 3'h0 == pht_windex & 8'hb7 == _GEN_14976 ? pht_0_183 : _GEN_2486; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15146 = 8'hb8 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2488 = 3'h0 == pht_windex & 8'hb8 == _GEN_14976 ? pht_0_184 : _GEN_2487; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15149 = 8'hb9 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2489 = 3'h0 == pht_windex & 8'hb9 == _GEN_14976 ? pht_0_185 : _GEN_2488; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15152 = 8'hba == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2490 = 3'h0 == pht_windex & 8'hba == _GEN_14976 ? pht_0_186 : _GEN_2489; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15155 = 8'hbb == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2491 = 3'h0 == pht_windex & 8'hbb == _GEN_14976 ? pht_0_187 : _GEN_2490; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15158 = 8'hbc == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2492 = 3'h0 == pht_windex & 8'hbc == _GEN_14976 ? pht_0_188 : _GEN_2491; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15161 = 8'hbd == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2493 = 3'h0 == pht_windex & 8'hbd == _GEN_14976 ? pht_0_189 : _GEN_2492; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15164 = 8'hbe == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2494 = 3'h0 == pht_windex & 8'hbe == _GEN_14976 ? pht_0_190 : _GEN_2493; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15167 = 8'hbf == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2495 = 3'h0 == pht_windex & 8'hbf == _GEN_14976 ? pht_0_191 : _GEN_2494; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15170 = 8'hc0 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2496 = 3'h0 == pht_windex & 8'hc0 == _GEN_14976 ? pht_0_192 : _GEN_2495; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15173 = 8'hc1 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2497 = 3'h0 == pht_windex & 8'hc1 == _GEN_14976 ? pht_0_193 : _GEN_2496; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15176 = 8'hc2 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2498 = 3'h0 == pht_windex & 8'hc2 == _GEN_14976 ? pht_0_194 : _GEN_2497; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15179 = 8'hc3 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2499 = 3'h0 == pht_windex & 8'hc3 == _GEN_14976 ? pht_0_195 : _GEN_2498; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15182 = 8'hc4 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2500 = 3'h0 == pht_windex & 8'hc4 == _GEN_14976 ? pht_0_196 : _GEN_2499; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15185 = 8'hc5 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2501 = 3'h0 == pht_windex & 8'hc5 == _GEN_14976 ? pht_0_197 : _GEN_2500; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15188 = 8'hc6 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2502 = 3'h0 == pht_windex & 8'hc6 == _GEN_14976 ? pht_0_198 : _GEN_2501; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15191 = 8'hc7 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2503 = 3'h0 == pht_windex & 8'hc7 == _GEN_14976 ? pht_0_199 : _GEN_2502; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15194 = 8'hc8 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2504 = 3'h0 == pht_windex & 8'hc8 == _GEN_14976 ? pht_0_200 : _GEN_2503; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15197 = 8'hc9 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2505 = 3'h0 == pht_windex & 8'hc9 == _GEN_14976 ? pht_0_201 : _GEN_2504; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15200 = 8'hca == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2506 = 3'h0 == pht_windex & 8'hca == _GEN_14976 ? pht_0_202 : _GEN_2505; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15203 = 8'hcb == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2507 = 3'h0 == pht_windex & 8'hcb == _GEN_14976 ? pht_0_203 : _GEN_2506; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15206 = 8'hcc == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2508 = 3'h0 == pht_windex & 8'hcc == _GEN_14976 ? pht_0_204 : _GEN_2507; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15209 = 8'hcd == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2509 = 3'h0 == pht_windex & 8'hcd == _GEN_14976 ? pht_0_205 : _GEN_2508; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15212 = 8'hce == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2510 = 3'h0 == pht_windex & 8'hce == _GEN_14976 ? pht_0_206 : _GEN_2509; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15215 = 8'hcf == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2511 = 3'h0 == pht_windex & 8'hcf == _GEN_14976 ? pht_0_207 : _GEN_2510; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15218 = 8'hd0 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2512 = 3'h0 == pht_windex & 8'hd0 == _GEN_14976 ? pht_0_208 : _GEN_2511; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15221 = 8'hd1 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2513 = 3'h0 == pht_windex & 8'hd1 == _GEN_14976 ? pht_0_209 : _GEN_2512; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15224 = 8'hd2 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2514 = 3'h0 == pht_windex & 8'hd2 == _GEN_14976 ? pht_0_210 : _GEN_2513; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15227 = 8'hd3 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2515 = 3'h0 == pht_windex & 8'hd3 == _GEN_14976 ? pht_0_211 : _GEN_2514; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15230 = 8'hd4 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2516 = 3'h0 == pht_windex & 8'hd4 == _GEN_14976 ? pht_0_212 : _GEN_2515; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15233 = 8'hd5 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2517 = 3'h0 == pht_windex & 8'hd5 == _GEN_14976 ? pht_0_213 : _GEN_2516; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15236 = 8'hd6 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2518 = 3'h0 == pht_windex & 8'hd6 == _GEN_14976 ? pht_0_214 : _GEN_2517; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15239 = 8'hd7 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2519 = 3'h0 == pht_windex & 8'hd7 == _GEN_14976 ? pht_0_215 : _GEN_2518; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15242 = 8'hd8 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2520 = 3'h0 == pht_windex & 8'hd8 == _GEN_14976 ? pht_0_216 : _GEN_2519; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15245 = 8'hd9 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2521 = 3'h0 == pht_windex & 8'hd9 == _GEN_14976 ? pht_0_217 : _GEN_2520; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15248 = 8'hda == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2522 = 3'h0 == pht_windex & 8'hda == _GEN_14976 ? pht_0_218 : _GEN_2521; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15251 = 8'hdb == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2523 = 3'h0 == pht_windex & 8'hdb == _GEN_14976 ? pht_0_219 : _GEN_2522; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15254 = 8'hdc == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2524 = 3'h0 == pht_windex & 8'hdc == _GEN_14976 ? pht_0_220 : _GEN_2523; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15257 = 8'hdd == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2525 = 3'h0 == pht_windex & 8'hdd == _GEN_14976 ? pht_0_221 : _GEN_2524; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15260 = 8'hde == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2526 = 3'h0 == pht_windex & 8'hde == _GEN_14976 ? pht_0_222 : _GEN_2525; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15263 = 8'hdf == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2527 = 3'h0 == pht_windex & 8'hdf == _GEN_14976 ? pht_0_223 : _GEN_2526; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15266 = 8'he0 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2528 = 3'h0 == pht_windex & 8'he0 == _GEN_14976 ? pht_0_224 : _GEN_2527; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15269 = 8'he1 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2529 = 3'h0 == pht_windex & 8'he1 == _GEN_14976 ? pht_0_225 : _GEN_2528; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15272 = 8'he2 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2530 = 3'h0 == pht_windex & 8'he2 == _GEN_14976 ? pht_0_226 : _GEN_2529; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15275 = 8'he3 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2531 = 3'h0 == pht_windex & 8'he3 == _GEN_14976 ? pht_0_227 : _GEN_2530; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15278 = 8'he4 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2532 = 3'h0 == pht_windex & 8'he4 == _GEN_14976 ? pht_0_228 : _GEN_2531; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15281 = 8'he5 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2533 = 3'h0 == pht_windex & 8'he5 == _GEN_14976 ? pht_0_229 : _GEN_2532; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15284 = 8'he6 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2534 = 3'h0 == pht_windex & 8'he6 == _GEN_14976 ? pht_0_230 : _GEN_2533; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15287 = 8'he7 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2535 = 3'h0 == pht_windex & 8'he7 == _GEN_14976 ? pht_0_231 : _GEN_2534; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15290 = 8'he8 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2536 = 3'h0 == pht_windex & 8'he8 == _GEN_14976 ? pht_0_232 : _GEN_2535; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15293 = 8'he9 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2537 = 3'h0 == pht_windex & 8'he9 == _GEN_14976 ? pht_0_233 : _GEN_2536; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15296 = 8'hea == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2538 = 3'h0 == pht_windex & 8'hea == _GEN_14976 ? pht_0_234 : _GEN_2537; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15299 = 8'heb == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2539 = 3'h0 == pht_windex & 8'heb == _GEN_14976 ? pht_0_235 : _GEN_2538; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15302 = 8'hec == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2540 = 3'h0 == pht_windex & 8'hec == _GEN_14976 ? pht_0_236 : _GEN_2539; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15305 = 8'hed == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2541 = 3'h0 == pht_windex & 8'hed == _GEN_14976 ? pht_0_237 : _GEN_2540; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15308 = 8'hee == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2542 = 3'h0 == pht_windex & 8'hee == _GEN_14976 ? pht_0_238 : _GEN_2541; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15311 = 8'hef == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2543 = 3'h0 == pht_windex & 8'hef == _GEN_14976 ? pht_0_239 : _GEN_2542; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15314 = 8'hf0 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2544 = 3'h0 == pht_windex & 8'hf0 == _GEN_14976 ? pht_0_240 : _GEN_2543; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15317 = 8'hf1 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2545 = 3'h0 == pht_windex & 8'hf1 == _GEN_14976 ? pht_0_241 : _GEN_2544; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15320 = 8'hf2 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2546 = 3'h0 == pht_windex & 8'hf2 == _GEN_14976 ? pht_0_242 : _GEN_2545; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15323 = 8'hf3 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2547 = 3'h0 == pht_windex & 8'hf3 == _GEN_14976 ? pht_0_243 : _GEN_2546; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15326 = 8'hf4 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2548 = 3'h0 == pht_windex & 8'hf4 == _GEN_14976 ? pht_0_244 : _GEN_2547; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15329 = 8'hf5 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2549 = 3'h0 == pht_windex & 8'hf5 == _GEN_14976 ? pht_0_245 : _GEN_2548; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15332 = 8'hf6 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2550 = 3'h0 == pht_windex & 8'hf6 == _GEN_14976 ? pht_0_246 : _GEN_2549; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15335 = 8'hf7 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2551 = 3'h0 == pht_windex & 8'hf7 == _GEN_14976 ? pht_0_247 : _GEN_2550; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15338 = 8'hf8 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2552 = 3'h0 == pht_windex & 8'hf8 == _GEN_14976 ? pht_0_248 : _GEN_2551; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15341 = 8'hf9 == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2553 = 3'h0 == pht_windex & 8'hf9 == _GEN_14976 ? pht_0_249 : _GEN_2552; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15344 = 8'hfa == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2554 = 3'h0 == pht_windex & 8'hfa == _GEN_14976 ? pht_0_250 : _GEN_2553; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15347 = 8'hfb == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2555 = 3'h0 == pht_windex & 8'hfb == _GEN_14976 ? pht_0_251 : _GEN_2554; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15350 = 8'hfc == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2556 = 3'h0 == pht_windex & 8'hfc == _GEN_14976 ? pht_0_252 : _GEN_2555; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15353 = 8'hfd == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2557 = 3'h0 == pht_windex & 8'hfd == _GEN_14976 ? pht_0_253 : _GEN_2556; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15356 = 8'hfe == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2558 = 3'h0 == pht_windex & 8'hfe == _GEN_14976 ? pht_0_254 : _GEN_2557; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15359 = 8'hff == _GEN_14976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2559 = 3'h0 == pht_windex & 8'hff == _GEN_14976 ? pht_0_255 : _GEN_2558; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15360 = 3'h1 == pht_windex; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_15361 = 6'h0 == pht_waddr; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2560 = 3'h1 == pht_windex & 6'h0 == pht_waddr ? pht_1_0 : _GEN_2559; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2561 = 3'h1 == pht_windex & 6'h1 == pht_waddr ? pht_1_1 : _GEN_2560; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2562 = 3'h1 == pht_windex & 6'h2 == pht_waddr ? pht_1_2 : _GEN_2561; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2563 = 3'h1 == pht_windex & 6'h3 == pht_waddr ? pht_1_3 : _GEN_2562; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2564 = 3'h1 == pht_windex & 6'h4 == pht_waddr ? pht_1_4 : _GEN_2563; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2565 = 3'h1 == pht_windex & 6'h5 == pht_waddr ? pht_1_5 : _GEN_2564; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2566 = 3'h1 == pht_windex & 6'h6 == pht_waddr ? pht_1_6 : _GEN_2565; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2567 = 3'h1 == pht_windex & 6'h7 == pht_waddr ? pht_1_7 : _GEN_2566; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2568 = 3'h1 == pht_windex & 6'h8 == pht_waddr ? pht_1_8 : _GEN_2567; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2569 = 3'h1 == pht_windex & 6'h9 == pht_waddr ? pht_1_9 : _GEN_2568; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2570 = 3'h1 == pht_windex & 6'ha == pht_waddr ? pht_1_10 : _GEN_2569; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2571 = 3'h1 == pht_windex & 6'hb == pht_waddr ? pht_1_11 : _GEN_2570; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2572 = 3'h1 == pht_windex & 6'hc == pht_waddr ? pht_1_12 : _GEN_2571; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2573 = 3'h1 == pht_windex & 6'hd == pht_waddr ? pht_1_13 : _GEN_2572; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2574 = 3'h1 == pht_windex & 6'he == pht_waddr ? pht_1_14 : _GEN_2573; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2575 = 3'h1 == pht_windex & 6'hf == pht_waddr ? pht_1_15 : _GEN_2574; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2576 = 3'h1 == pht_windex & 6'h10 == pht_waddr ? pht_1_16 : _GEN_2575; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2577 = 3'h1 == pht_windex & 6'h11 == pht_waddr ? pht_1_17 : _GEN_2576; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2578 = 3'h1 == pht_windex & 6'h12 == pht_waddr ? pht_1_18 : _GEN_2577; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2579 = 3'h1 == pht_windex & 6'h13 == pht_waddr ? pht_1_19 : _GEN_2578; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2580 = 3'h1 == pht_windex & 6'h14 == pht_waddr ? pht_1_20 : _GEN_2579; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2581 = 3'h1 == pht_windex & 6'h15 == pht_waddr ? pht_1_21 : _GEN_2580; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2582 = 3'h1 == pht_windex & 6'h16 == pht_waddr ? pht_1_22 : _GEN_2581; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2583 = 3'h1 == pht_windex & 6'h17 == pht_waddr ? pht_1_23 : _GEN_2582; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2584 = 3'h1 == pht_windex & 6'h18 == pht_waddr ? pht_1_24 : _GEN_2583; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2585 = 3'h1 == pht_windex & 6'h19 == pht_waddr ? pht_1_25 : _GEN_2584; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2586 = 3'h1 == pht_windex & 6'h1a == pht_waddr ? pht_1_26 : _GEN_2585; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2587 = 3'h1 == pht_windex & 6'h1b == pht_waddr ? pht_1_27 : _GEN_2586; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2588 = 3'h1 == pht_windex & 6'h1c == pht_waddr ? pht_1_28 : _GEN_2587; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2589 = 3'h1 == pht_windex & 6'h1d == pht_waddr ? pht_1_29 : _GEN_2588; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2590 = 3'h1 == pht_windex & 6'h1e == pht_waddr ? pht_1_30 : _GEN_2589; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2591 = 3'h1 == pht_windex & 6'h1f == pht_waddr ? pht_1_31 : _GEN_2590; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2592 = 3'h1 == pht_windex & 6'h20 == pht_waddr ? pht_1_32 : _GEN_2591; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2593 = 3'h1 == pht_windex & 6'h21 == pht_waddr ? pht_1_33 : _GEN_2592; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2594 = 3'h1 == pht_windex & 6'h22 == pht_waddr ? pht_1_34 : _GEN_2593; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2595 = 3'h1 == pht_windex & 6'h23 == pht_waddr ? pht_1_35 : _GEN_2594; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2596 = 3'h1 == pht_windex & 6'h24 == pht_waddr ? pht_1_36 : _GEN_2595; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2597 = 3'h1 == pht_windex & 6'h25 == pht_waddr ? pht_1_37 : _GEN_2596; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2598 = 3'h1 == pht_windex & 6'h26 == pht_waddr ? pht_1_38 : _GEN_2597; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2599 = 3'h1 == pht_windex & 6'h27 == pht_waddr ? pht_1_39 : _GEN_2598; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2600 = 3'h1 == pht_windex & 6'h28 == pht_waddr ? pht_1_40 : _GEN_2599; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2601 = 3'h1 == pht_windex & 6'h29 == pht_waddr ? pht_1_41 : _GEN_2600; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2602 = 3'h1 == pht_windex & 6'h2a == pht_waddr ? pht_1_42 : _GEN_2601; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2603 = 3'h1 == pht_windex & 6'h2b == pht_waddr ? pht_1_43 : _GEN_2602; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2604 = 3'h1 == pht_windex & 6'h2c == pht_waddr ? pht_1_44 : _GEN_2603; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2605 = 3'h1 == pht_windex & 6'h2d == pht_waddr ? pht_1_45 : _GEN_2604; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2606 = 3'h1 == pht_windex & 6'h2e == pht_waddr ? pht_1_46 : _GEN_2605; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2607 = 3'h1 == pht_windex & 6'h2f == pht_waddr ? pht_1_47 : _GEN_2606; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2608 = 3'h1 == pht_windex & 6'h30 == pht_waddr ? pht_1_48 : _GEN_2607; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2609 = 3'h1 == pht_windex & 6'h31 == pht_waddr ? pht_1_49 : _GEN_2608; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2610 = 3'h1 == pht_windex & 6'h32 == pht_waddr ? pht_1_50 : _GEN_2609; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2611 = 3'h1 == pht_windex & 6'h33 == pht_waddr ? pht_1_51 : _GEN_2610; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2612 = 3'h1 == pht_windex & 6'h34 == pht_waddr ? pht_1_52 : _GEN_2611; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2613 = 3'h1 == pht_windex & 6'h35 == pht_waddr ? pht_1_53 : _GEN_2612; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2614 = 3'h1 == pht_windex & 6'h36 == pht_waddr ? pht_1_54 : _GEN_2613; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2615 = 3'h1 == pht_windex & 6'h37 == pht_waddr ? pht_1_55 : _GEN_2614; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2616 = 3'h1 == pht_windex & 6'h38 == pht_waddr ? pht_1_56 : _GEN_2615; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2617 = 3'h1 == pht_windex & 6'h39 == pht_waddr ? pht_1_57 : _GEN_2616; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2618 = 3'h1 == pht_windex & 6'h3a == pht_waddr ? pht_1_58 : _GEN_2617; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2619 = 3'h1 == pht_windex & 6'h3b == pht_waddr ? pht_1_59 : _GEN_2618; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2620 = 3'h1 == pht_windex & 6'h3c == pht_waddr ? pht_1_60 : _GEN_2619; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2621 = 3'h1 == pht_windex & 6'h3d == pht_waddr ? pht_1_61 : _GEN_2620; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2622 = 3'h1 == pht_windex & 6'h3e == pht_waddr ? pht_1_62 : _GEN_2621; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2623 = 3'h1 == pht_windex & 6'h3f == pht_waddr ? pht_1_63 : _GEN_2622; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2624 = 3'h1 == pht_windex & 7'h40 == _GEN_14784 ? pht_1_64 : _GEN_2623; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2625 = 3'h1 == pht_windex & 7'h41 == _GEN_14784 ? pht_1_65 : _GEN_2624; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2626 = 3'h1 == pht_windex & 7'h42 == _GEN_14784 ? pht_1_66 : _GEN_2625; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2627 = 3'h1 == pht_windex & 7'h43 == _GEN_14784 ? pht_1_67 : _GEN_2626; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2628 = 3'h1 == pht_windex & 7'h44 == _GEN_14784 ? pht_1_68 : _GEN_2627; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2629 = 3'h1 == pht_windex & 7'h45 == _GEN_14784 ? pht_1_69 : _GEN_2628; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2630 = 3'h1 == pht_windex & 7'h46 == _GEN_14784 ? pht_1_70 : _GEN_2629; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2631 = 3'h1 == pht_windex & 7'h47 == _GEN_14784 ? pht_1_71 : _GEN_2630; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2632 = 3'h1 == pht_windex & 7'h48 == _GEN_14784 ? pht_1_72 : _GEN_2631; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2633 = 3'h1 == pht_windex & 7'h49 == _GEN_14784 ? pht_1_73 : _GEN_2632; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2634 = 3'h1 == pht_windex & 7'h4a == _GEN_14784 ? pht_1_74 : _GEN_2633; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2635 = 3'h1 == pht_windex & 7'h4b == _GEN_14784 ? pht_1_75 : _GEN_2634; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2636 = 3'h1 == pht_windex & 7'h4c == _GEN_14784 ? pht_1_76 : _GEN_2635; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2637 = 3'h1 == pht_windex & 7'h4d == _GEN_14784 ? pht_1_77 : _GEN_2636; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2638 = 3'h1 == pht_windex & 7'h4e == _GEN_14784 ? pht_1_78 : _GEN_2637; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2639 = 3'h1 == pht_windex & 7'h4f == _GEN_14784 ? pht_1_79 : _GEN_2638; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2640 = 3'h1 == pht_windex & 7'h50 == _GEN_14784 ? pht_1_80 : _GEN_2639; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2641 = 3'h1 == pht_windex & 7'h51 == _GEN_14784 ? pht_1_81 : _GEN_2640; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2642 = 3'h1 == pht_windex & 7'h52 == _GEN_14784 ? pht_1_82 : _GEN_2641; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2643 = 3'h1 == pht_windex & 7'h53 == _GEN_14784 ? pht_1_83 : _GEN_2642; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2644 = 3'h1 == pht_windex & 7'h54 == _GEN_14784 ? pht_1_84 : _GEN_2643; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2645 = 3'h1 == pht_windex & 7'h55 == _GEN_14784 ? pht_1_85 : _GEN_2644; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2646 = 3'h1 == pht_windex & 7'h56 == _GEN_14784 ? pht_1_86 : _GEN_2645; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2647 = 3'h1 == pht_windex & 7'h57 == _GEN_14784 ? pht_1_87 : _GEN_2646; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2648 = 3'h1 == pht_windex & 7'h58 == _GEN_14784 ? pht_1_88 : _GEN_2647; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2649 = 3'h1 == pht_windex & 7'h59 == _GEN_14784 ? pht_1_89 : _GEN_2648; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2650 = 3'h1 == pht_windex & 7'h5a == _GEN_14784 ? pht_1_90 : _GEN_2649; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2651 = 3'h1 == pht_windex & 7'h5b == _GEN_14784 ? pht_1_91 : _GEN_2650; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2652 = 3'h1 == pht_windex & 7'h5c == _GEN_14784 ? pht_1_92 : _GEN_2651; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2653 = 3'h1 == pht_windex & 7'h5d == _GEN_14784 ? pht_1_93 : _GEN_2652; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2654 = 3'h1 == pht_windex & 7'h5e == _GEN_14784 ? pht_1_94 : _GEN_2653; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2655 = 3'h1 == pht_windex & 7'h5f == _GEN_14784 ? pht_1_95 : _GEN_2654; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2656 = 3'h1 == pht_windex & 7'h60 == _GEN_14784 ? pht_1_96 : _GEN_2655; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2657 = 3'h1 == pht_windex & 7'h61 == _GEN_14784 ? pht_1_97 : _GEN_2656; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2658 = 3'h1 == pht_windex & 7'h62 == _GEN_14784 ? pht_1_98 : _GEN_2657; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2659 = 3'h1 == pht_windex & 7'h63 == _GEN_14784 ? pht_1_99 : _GEN_2658; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2660 = 3'h1 == pht_windex & 7'h64 == _GEN_14784 ? pht_1_100 : _GEN_2659; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2661 = 3'h1 == pht_windex & 7'h65 == _GEN_14784 ? pht_1_101 : _GEN_2660; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2662 = 3'h1 == pht_windex & 7'h66 == _GEN_14784 ? pht_1_102 : _GEN_2661; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2663 = 3'h1 == pht_windex & 7'h67 == _GEN_14784 ? pht_1_103 : _GEN_2662; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2664 = 3'h1 == pht_windex & 7'h68 == _GEN_14784 ? pht_1_104 : _GEN_2663; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2665 = 3'h1 == pht_windex & 7'h69 == _GEN_14784 ? pht_1_105 : _GEN_2664; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2666 = 3'h1 == pht_windex & 7'h6a == _GEN_14784 ? pht_1_106 : _GEN_2665; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2667 = 3'h1 == pht_windex & 7'h6b == _GEN_14784 ? pht_1_107 : _GEN_2666; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2668 = 3'h1 == pht_windex & 7'h6c == _GEN_14784 ? pht_1_108 : _GEN_2667; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2669 = 3'h1 == pht_windex & 7'h6d == _GEN_14784 ? pht_1_109 : _GEN_2668; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2670 = 3'h1 == pht_windex & 7'h6e == _GEN_14784 ? pht_1_110 : _GEN_2669; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2671 = 3'h1 == pht_windex & 7'h6f == _GEN_14784 ? pht_1_111 : _GEN_2670; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2672 = 3'h1 == pht_windex & 7'h70 == _GEN_14784 ? pht_1_112 : _GEN_2671; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2673 = 3'h1 == pht_windex & 7'h71 == _GEN_14784 ? pht_1_113 : _GEN_2672; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2674 = 3'h1 == pht_windex & 7'h72 == _GEN_14784 ? pht_1_114 : _GEN_2673; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2675 = 3'h1 == pht_windex & 7'h73 == _GEN_14784 ? pht_1_115 : _GEN_2674; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2676 = 3'h1 == pht_windex & 7'h74 == _GEN_14784 ? pht_1_116 : _GEN_2675; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2677 = 3'h1 == pht_windex & 7'h75 == _GEN_14784 ? pht_1_117 : _GEN_2676; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2678 = 3'h1 == pht_windex & 7'h76 == _GEN_14784 ? pht_1_118 : _GEN_2677; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2679 = 3'h1 == pht_windex & 7'h77 == _GEN_14784 ? pht_1_119 : _GEN_2678; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2680 = 3'h1 == pht_windex & 7'h78 == _GEN_14784 ? pht_1_120 : _GEN_2679; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2681 = 3'h1 == pht_windex & 7'h79 == _GEN_14784 ? pht_1_121 : _GEN_2680; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2682 = 3'h1 == pht_windex & 7'h7a == _GEN_14784 ? pht_1_122 : _GEN_2681; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2683 = 3'h1 == pht_windex & 7'h7b == _GEN_14784 ? pht_1_123 : _GEN_2682; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2684 = 3'h1 == pht_windex & 7'h7c == _GEN_14784 ? pht_1_124 : _GEN_2683; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2685 = 3'h1 == pht_windex & 7'h7d == _GEN_14784 ? pht_1_125 : _GEN_2684; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2686 = 3'h1 == pht_windex & 7'h7e == _GEN_14784 ? pht_1_126 : _GEN_2685; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2687 = 3'h1 == pht_windex & 7'h7f == _GEN_14784 ? pht_1_127 : _GEN_2686; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2688 = 3'h1 == pht_windex & 8'h80 == _GEN_14976 ? pht_1_128 : _GEN_2687; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2689 = 3'h1 == pht_windex & 8'h81 == _GEN_14976 ? pht_1_129 : _GEN_2688; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2690 = 3'h1 == pht_windex & 8'h82 == _GEN_14976 ? pht_1_130 : _GEN_2689; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2691 = 3'h1 == pht_windex & 8'h83 == _GEN_14976 ? pht_1_131 : _GEN_2690; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2692 = 3'h1 == pht_windex & 8'h84 == _GEN_14976 ? pht_1_132 : _GEN_2691; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2693 = 3'h1 == pht_windex & 8'h85 == _GEN_14976 ? pht_1_133 : _GEN_2692; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2694 = 3'h1 == pht_windex & 8'h86 == _GEN_14976 ? pht_1_134 : _GEN_2693; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2695 = 3'h1 == pht_windex & 8'h87 == _GEN_14976 ? pht_1_135 : _GEN_2694; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2696 = 3'h1 == pht_windex & 8'h88 == _GEN_14976 ? pht_1_136 : _GEN_2695; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2697 = 3'h1 == pht_windex & 8'h89 == _GEN_14976 ? pht_1_137 : _GEN_2696; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2698 = 3'h1 == pht_windex & 8'h8a == _GEN_14976 ? pht_1_138 : _GEN_2697; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2699 = 3'h1 == pht_windex & 8'h8b == _GEN_14976 ? pht_1_139 : _GEN_2698; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2700 = 3'h1 == pht_windex & 8'h8c == _GEN_14976 ? pht_1_140 : _GEN_2699; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2701 = 3'h1 == pht_windex & 8'h8d == _GEN_14976 ? pht_1_141 : _GEN_2700; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2702 = 3'h1 == pht_windex & 8'h8e == _GEN_14976 ? pht_1_142 : _GEN_2701; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2703 = 3'h1 == pht_windex & 8'h8f == _GEN_14976 ? pht_1_143 : _GEN_2702; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2704 = 3'h1 == pht_windex & 8'h90 == _GEN_14976 ? pht_1_144 : _GEN_2703; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2705 = 3'h1 == pht_windex & 8'h91 == _GEN_14976 ? pht_1_145 : _GEN_2704; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2706 = 3'h1 == pht_windex & 8'h92 == _GEN_14976 ? pht_1_146 : _GEN_2705; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2707 = 3'h1 == pht_windex & 8'h93 == _GEN_14976 ? pht_1_147 : _GEN_2706; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2708 = 3'h1 == pht_windex & 8'h94 == _GEN_14976 ? pht_1_148 : _GEN_2707; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2709 = 3'h1 == pht_windex & 8'h95 == _GEN_14976 ? pht_1_149 : _GEN_2708; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2710 = 3'h1 == pht_windex & 8'h96 == _GEN_14976 ? pht_1_150 : _GEN_2709; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2711 = 3'h1 == pht_windex & 8'h97 == _GEN_14976 ? pht_1_151 : _GEN_2710; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2712 = 3'h1 == pht_windex & 8'h98 == _GEN_14976 ? pht_1_152 : _GEN_2711; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2713 = 3'h1 == pht_windex & 8'h99 == _GEN_14976 ? pht_1_153 : _GEN_2712; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2714 = 3'h1 == pht_windex & 8'h9a == _GEN_14976 ? pht_1_154 : _GEN_2713; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2715 = 3'h1 == pht_windex & 8'h9b == _GEN_14976 ? pht_1_155 : _GEN_2714; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2716 = 3'h1 == pht_windex & 8'h9c == _GEN_14976 ? pht_1_156 : _GEN_2715; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2717 = 3'h1 == pht_windex & 8'h9d == _GEN_14976 ? pht_1_157 : _GEN_2716; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2718 = 3'h1 == pht_windex & 8'h9e == _GEN_14976 ? pht_1_158 : _GEN_2717; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2719 = 3'h1 == pht_windex & 8'h9f == _GEN_14976 ? pht_1_159 : _GEN_2718; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2720 = 3'h1 == pht_windex & 8'ha0 == _GEN_14976 ? pht_1_160 : _GEN_2719; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2721 = 3'h1 == pht_windex & 8'ha1 == _GEN_14976 ? pht_1_161 : _GEN_2720; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2722 = 3'h1 == pht_windex & 8'ha2 == _GEN_14976 ? pht_1_162 : _GEN_2721; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2723 = 3'h1 == pht_windex & 8'ha3 == _GEN_14976 ? pht_1_163 : _GEN_2722; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2724 = 3'h1 == pht_windex & 8'ha4 == _GEN_14976 ? pht_1_164 : _GEN_2723; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2725 = 3'h1 == pht_windex & 8'ha5 == _GEN_14976 ? pht_1_165 : _GEN_2724; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2726 = 3'h1 == pht_windex & 8'ha6 == _GEN_14976 ? pht_1_166 : _GEN_2725; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2727 = 3'h1 == pht_windex & 8'ha7 == _GEN_14976 ? pht_1_167 : _GEN_2726; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2728 = 3'h1 == pht_windex & 8'ha8 == _GEN_14976 ? pht_1_168 : _GEN_2727; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2729 = 3'h1 == pht_windex & 8'ha9 == _GEN_14976 ? pht_1_169 : _GEN_2728; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2730 = 3'h1 == pht_windex & 8'haa == _GEN_14976 ? pht_1_170 : _GEN_2729; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2731 = 3'h1 == pht_windex & 8'hab == _GEN_14976 ? pht_1_171 : _GEN_2730; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2732 = 3'h1 == pht_windex & 8'hac == _GEN_14976 ? pht_1_172 : _GEN_2731; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2733 = 3'h1 == pht_windex & 8'had == _GEN_14976 ? pht_1_173 : _GEN_2732; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2734 = 3'h1 == pht_windex & 8'hae == _GEN_14976 ? pht_1_174 : _GEN_2733; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2735 = 3'h1 == pht_windex & 8'haf == _GEN_14976 ? pht_1_175 : _GEN_2734; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2736 = 3'h1 == pht_windex & 8'hb0 == _GEN_14976 ? pht_1_176 : _GEN_2735; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2737 = 3'h1 == pht_windex & 8'hb1 == _GEN_14976 ? pht_1_177 : _GEN_2736; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2738 = 3'h1 == pht_windex & 8'hb2 == _GEN_14976 ? pht_1_178 : _GEN_2737; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2739 = 3'h1 == pht_windex & 8'hb3 == _GEN_14976 ? pht_1_179 : _GEN_2738; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2740 = 3'h1 == pht_windex & 8'hb4 == _GEN_14976 ? pht_1_180 : _GEN_2739; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2741 = 3'h1 == pht_windex & 8'hb5 == _GEN_14976 ? pht_1_181 : _GEN_2740; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2742 = 3'h1 == pht_windex & 8'hb6 == _GEN_14976 ? pht_1_182 : _GEN_2741; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2743 = 3'h1 == pht_windex & 8'hb7 == _GEN_14976 ? pht_1_183 : _GEN_2742; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2744 = 3'h1 == pht_windex & 8'hb8 == _GEN_14976 ? pht_1_184 : _GEN_2743; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2745 = 3'h1 == pht_windex & 8'hb9 == _GEN_14976 ? pht_1_185 : _GEN_2744; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2746 = 3'h1 == pht_windex & 8'hba == _GEN_14976 ? pht_1_186 : _GEN_2745; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2747 = 3'h1 == pht_windex & 8'hbb == _GEN_14976 ? pht_1_187 : _GEN_2746; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2748 = 3'h1 == pht_windex & 8'hbc == _GEN_14976 ? pht_1_188 : _GEN_2747; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2749 = 3'h1 == pht_windex & 8'hbd == _GEN_14976 ? pht_1_189 : _GEN_2748; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2750 = 3'h1 == pht_windex & 8'hbe == _GEN_14976 ? pht_1_190 : _GEN_2749; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2751 = 3'h1 == pht_windex & 8'hbf == _GEN_14976 ? pht_1_191 : _GEN_2750; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2752 = 3'h1 == pht_windex & 8'hc0 == _GEN_14976 ? pht_1_192 : _GEN_2751; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2753 = 3'h1 == pht_windex & 8'hc1 == _GEN_14976 ? pht_1_193 : _GEN_2752; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2754 = 3'h1 == pht_windex & 8'hc2 == _GEN_14976 ? pht_1_194 : _GEN_2753; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2755 = 3'h1 == pht_windex & 8'hc3 == _GEN_14976 ? pht_1_195 : _GEN_2754; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2756 = 3'h1 == pht_windex & 8'hc4 == _GEN_14976 ? pht_1_196 : _GEN_2755; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2757 = 3'h1 == pht_windex & 8'hc5 == _GEN_14976 ? pht_1_197 : _GEN_2756; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2758 = 3'h1 == pht_windex & 8'hc6 == _GEN_14976 ? pht_1_198 : _GEN_2757; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2759 = 3'h1 == pht_windex & 8'hc7 == _GEN_14976 ? pht_1_199 : _GEN_2758; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2760 = 3'h1 == pht_windex & 8'hc8 == _GEN_14976 ? pht_1_200 : _GEN_2759; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2761 = 3'h1 == pht_windex & 8'hc9 == _GEN_14976 ? pht_1_201 : _GEN_2760; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2762 = 3'h1 == pht_windex & 8'hca == _GEN_14976 ? pht_1_202 : _GEN_2761; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2763 = 3'h1 == pht_windex & 8'hcb == _GEN_14976 ? pht_1_203 : _GEN_2762; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2764 = 3'h1 == pht_windex & 8'hcc == _GEN_14976 ? pht_1_204 : _GEN_2763; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2765 = 3'h1 == pht_windex & 8'hcd == _GEN_14976 ? pht_1_205 : _GEN_2764; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2766 = 3'h1 == pht_windex & 8'hce == _GEN_14976 ? pht_1_206 : _GEN_2765; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2767 = 3'h1 == pht_windex & 8'hcf == _GEN_14976 ? pht_1_207 : _GEN_2766; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2768 = 3'h1 == pht_windex & 8'hd0 == _GEN_14976 ? pht_1_208 : _GEN_2767; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2769 = 3'h1 == pht_windex & 8'hd1 == _GEN_14976 ? pht_1_209 : _GEN_2768; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2770 = 3'h1 == pht_windex & 8'hd2 == _GEN_14976 ? pht_1_210 : _GEN_2769; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2771 = 3'h1 == pht_windex & 8'hd3 == _GEN_14976 ? pht_1_211 : _GEN_2770; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2772 = 3'h1 == pht_windex & 8'hd4 == _GEN_14976 ? pht_1_212 : _GEN_2771; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2773 = 3'h1 == pht_windex & 8'hd5 == _GEN_14976 ? pht_1_213 : _GEN_2772; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2774 = 3'h1 == pht_windex & 8'hd6 == _GEN_14976 ? pht_1_214 : _GEN_2773; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2775 = 3'h1 == pht_windex & 8'hd7 == _GEN_14976 ? pht_1_215 : _GEN_2774; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2776 = 3'h1 == pht_windex & 8'hd8 == _GEN_14976 ? pht_1_216 : _GEN_2775; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2777 = 3'h1 == pht_windex & 8'hd9 == _GEN_14976 ? pht_1_217 : _GEN_2776; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2778 = 3'h1 == pht_windex & 8'hda == _GEN_14976 ? pht_1_218 : _GEN_2777; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2779 = 3'h1 == pht_windex & 8'hdb == _GEN_14976 ? pht_1_219 : _GEN_2778; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2780 = 3'h1 == pht_windex & 8'hdc == _GEN_14976 ? pht_1_220 : _GEN_2779; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2781 = 3'h1 == pht_windex & 8'hdd == _GEN_14976 ? pht_1_221 : _GEN_2780; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2782 = 3'h1 == pht_windex & 8'hde == _GEN_14976 ? pht_1_222 : _GEN_2781; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2783 = 3'h1 == pht_windex & 8'hdf == _GEN_14976 ? pht_1_223 : _GEN_2782; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2784 = 3'h1 == pht_windex & 8'he0 == _GEN_14976 ? pht_1_224 : _GEN_2783; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2785 = 3'h1 == pht_windex & 8'he1 == _GEN_14976 ? pht_1_225 : _GEN_2784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2786 = 3'h1 == pht_windex & 8'he2 == _GEN_14976 ? pht_1_226 : _GEN_2785; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2787 = 3'h1 == pht_windex & 8'he3 == _GEN_14976 ? pht_1_227 : _GEN_2786; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2788 = 3'h1 == pht_windex & 8'he4 == _GEN_14976 ? pht_1_228 : _GEN_2787; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2789 = 3'h1 == pht_windex & 8'he5 == _GEN_14976 ? pht_1_229 : _GEN_2788; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2790 = 3'h1 == pht_windex & 8'he6 == _GEN_14976 ? pht_1_230 : _GEN_2789; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2791 = 3'h1 == pht_windex & 8'he7 == _GEN_14976 ? pht_1_231 : _GEN_2790; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2792 = 3'h1 == pht_windex & 8'he8 == _GEN_14976 ? pht_1_232 : _GEN_2791; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2793 = 3'h1 == pht_windex & 8'he9 == _GEN_14976 ? pht_1_233 : _GEN_2792; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2794 = 3'h1 == pht_windex & 8'hea == _GEN_14976 ? pht_1_234 : _GEN_2793; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2795 = 3'h1 == pht_windex & 8'heb == _GEN_14976 ? pht_1_235 : _GEN_2794; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2796 = 3'h1 == pht_windex & 8'hec == _GEN_14976 ? pht_1_236 : _GEN_2795; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2797 = 3'h1 == pht_windex & 8'hed == _GEN_14976 ? pht_1_237 : _GEN_2796; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2798 = 3'h1 == pht_windex & 8'hee == _GEN_14976 ? pht_1_238 : _GEN_2797; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2799 = 3'h1 == pht_windex & 8'hef == _GEN_14976 ? pht_1_239 : _GEN_2798; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2800 = 3'h1 == pht_windex & 8'hf0 == _GEN_14976 ? pht_1_240 : _GEN_2799; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2801 = 3'h1 == pht_windex & 8'hf1 == _GEN_14976 ? pht_1_241 : _GEN_2800; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2802 = 3'h1 == pht_windex & 8'hf2 == _GEN_14976 ? pht_1_242 : _GEN_2801; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2803 = 3'h1 == pht_windex & 8'hf3 == _GEN_14976 ? pht_1_243 : _GEN_2802; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2804 = 3'h1 == pht_windex & 8'hf4 == _GEN_14976 ? pht_1_244 : _GEN_2803; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2805 = 3'h1 == pht_windex & 8'hf5 == _GEN_14976 ? pht_1_245 : _GEN_2804; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2806 = 3'h1 == pht_windex & 8'hf6 == _GEN_14976 ? pht_1_246 : _GEN_2805; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2807 = 3'h1 == pht_windex & 8'hf7 == _GEN_14976 ? pht_1_247 : _GEN_2806; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2808 = 3'h1 == pht_windex & 8'hf8 == _GEN_14976 ? pht_1_248 : _GEN_2807; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2809 = 3'h1 == pht_windex & 8'hf9 == _GEN_14976 ? pht_1_249 : _GEN_2808; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2810 = 3'h1 == pht_windex & 8'hfa == _GEN_14976 ? pht_1_250 : _GEN_2809; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2811 = 3'h1 == pht_windex & 8'hfb == _GEN_14976 ? pht_1_251 : _GEN_2810; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2812 = 3'h1 == pht_windex & 8'hfc == _GEN_14976 ? pht_1_252 : _GEN_2811; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2813 = 3'h1 == pht_windex & 8'hfd == _GEN_14976 ? pht_1_253 : _GEN_2812; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2814 = 3'h1 == pht_windex & 8'hfe == _GEN_14976 ? pht_1_254 : _GEN_2813; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2815 = 3'h1 == pht_windex & 8'hff == _GEN_14976 ? pht_1_255 : _GEN_2814; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_16064 = 3'h2 == pht_windex; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2816 = 3'h2 == pht_windex & 6'h0 == pht_waddr ? pht_2_0 : _GEN_2815; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2817 = 3'h2 == pht_windex & 6'h1 == pht_waddr ? pht_2_1 : _GEN_2816; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2818 = 3'h2 == pht_windex & 6'h2 == pht_waddr ? pht_2_2 : _GEN_2817; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2819 = 3'h2 == pht_windex & 6'h3 == pht_waddr ? pht_2_3 : _GEN_2818; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2820 = 3'h2 == pht_windex & 6'h4 == pht_waddr ? pht_2_4 : _GEN_2819; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2821 = 3'h2 == pht_windex & 6'h5 == pht_waddr ? pht_2_5 : _GEN_2820; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2822 = 3'h2 == pht_windex & 6'h6 == pht_waddr ? pht_2_6 : _GEN_2821; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2823 = 3'h2 == pht_windex & 6'h7 == pht_waddr ? pht_2_7 : _GEN_2822; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2824 = 3'h2 == pht_windex & 6'h8 == pht_waddr ? pht_2_8 : _GEN_2823; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2825 = 3'h2 == pht_windex & 6'h9 == pht_waddr ? pht_2_9 : _GEN_2824; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2826 = 3'h2 == pht_windex & 6'ha == pht_waddr ? pht_2_10 : _GEN_2825; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2827 = 3'h2 == pht_windex & 6'hb == pht_waddr ? pht_2_11 : _GEN_2826; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2828 = 3'h2 == pht_windex & 6'hc == pht_waddr ? pht_2_12 : _GEN_2827; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2829 = 3'h2 == pht_windex & 6'hd == pht_waddr ? pht_2_13 : _GEN_2828; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2830 = 3'h2 == pht_windex & 6'he == pht_waddr ? pht_2_14 : _GEN_2829; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2831 = 3'h2 == pht_windex & 6'hf == pht_waddr ? pht_2_15 : _GEN_2830; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2832 = 3'h2 == pht_windex & 6'h10 == pht_waddr ? pht_2_16 : _GEN_2831; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2833 = 3'h2 == pht_windex & 6'h11 == pht_waddr ? pht_2_17 : _GEN_2832; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2834 = 3'h2 == pht_windex & 6'h12 == pht_waddr ? pht_2_18 : _GEN_2833; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2835 = 3'h2 == pht_windex & 6'h13 == pht_waddr ? pht_2_19 : _GEN_2834; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2836 = 3'h2 == pht_windex & 6'h14 == pht_waddr ? pht_2_20 : _GEN_2835; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2837 = 3'h2 == pht_windex & 6'h15 == pht_waddr ? pht_2_21 : _GEN_2836; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2838 = 3'h2 == pht_windex & 6'h16 == pht_waddr ? pht_2_22 : _GEN_2837; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2839 = 3'h2 == pht_windex & 6'h17 == pht_waddr ? pht_2_23 : _GEN_2838; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2840 = 3'h2 == pht_windex & 6'h18 == pht_waddr ? pht_2_24 : _GEN_2839; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2841 = 3'h2 == pht_windex & 6'h19 == pht_waddr ? pht_2_25 : _GEN_2840; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2842 = 3'h2 == pht_windex & 6'h1a == pht_waddr ? pht_2_26 : _GEN_2841; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2843 = 3'h2 == pht_windex & 6'h1b == pht_waddr ? pht_2_27 : _GEN_2842; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2844 = 3'h2 == pht_windex & 6'h1c == pht_waddr ? pht_2_28 : _GEN_2843; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2845 = 3'h2 == pht_windex & 6'h1d == pht_waddr ? pht_2_29 : _GEN_2844; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2846 = 3'h2 == pht_windex & 6'h1e == pht_waddr ? pht_2_30 : _GEN_2845; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2847 = 3'h2 == pht_windex & 6'h1f == pht_waddr ? pht_2_31 : _GEN_2846; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2848 = 3'h2 == pht_windex & 6'h20 == pht_waddr ? pht_2_32 : _GEN_2847; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2849 = 3'h2 == pht_windex & 6'h21 == pht_waddr ? pht_2_33 : _GEN_2848; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2850 = 3'h2 == pht_windex & 6'h22 == pht_waddr ? pht_2_34 : _GEN_2849; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2851 = 3'h2 == pht_windex & 6'h23 == pht_waddr ? pht_2_35 : _GEN_2850; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2852 = 3'h2 == pht_windex & 6'h24 == pht_waddr ? pht_2_36 : _GEN_2851; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2853 = 3'h2 == pht_windex & 6'h25 == pht_waddr ? pht_2_37 : _GEN_2852; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2854 = 3'h2 == pht_windex & 6'h26 == pht_waddr ? pht_2_38 : _GEN_2853; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2855 = 3'h2 == pht_windex & 6'h27 == pht_waddr ? pht_2_39 : _GEN_2854; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2856 = 3'h2 == pht_windex & 6'h28 == pht_waddr ? pht_2_40 : _GEN_2855; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2857 = 3'h2 == pht_windex & 6'h29 == pht_waddr ? pht_2_41 : _GEN_2856; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2858 = 3'h2 == pht_windex & 6'h2a == pht_waddr ? pht_2_42 : _GEN_2857; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2859 = 3'h2 == pht_windex & 6'h2b == pht_waddr ? pht_2_43 : _GEN_2858; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2860 = 3'h2 == pht_windex & 6'h2c == pht_waddr ? pht_2_44 : _GEN_2859; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2861 = 3'h2 == pht_windex & 6'h2d == pht_waddr ? pht_2_45 : _GEN_2860; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2862 = 3'h2 == pht_windex & 6'h2e == pht_waddr ? pht_2_46 : _GEN_2861; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2863 = 3'h2 == pht_windex & 6'h2f == pht_waddr ? pht_2_47 : _GEN_2862; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2864 = 3'h2 == pht_windex & 6'h30 == pht_waddr ? pht_2_48 : _GEN_2863; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2865 = 3'h2 == pht_windex & 6'h31 == pht_waddr ? pht_2_49 : _GEN_2864; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2866 = 3'h2 == pht_windex & 6'h32 == pht_waddr ? pht_2_50 : _GEN_2865; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2867 = 3'h2 == pht_windex & 6'h33 == pht_waddr ? pht_2_51 : _GEN_2866; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2868 = 3'h2 == pht_windex & 6'h34 == pht_waddr ? pht_2_52 : _GEN_2867; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2869 = 3'h2 == pht_windex & 6'h35 == pht_waddr ? pht_2_53 : _GEN_2868; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2870 = 3'h2 == pht_windex & 6'h36 == pht_waddr ? pht_2_54 : _GEN_2869; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2871 = 3'h2 == pht_windex & 6'h37 == pht_waddr ? pht_2_55 : _GEN_2870; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2872 = 3'h2 == pht_windex & 6'h38 == pht_waddr ? pht_2_56 : _GEN_2871; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2873 = 3'h2 == pht_windex & 6'h39 == pht_waddr ? pht_2_57 : _GEN_2872; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2874 = 3'h2 == pht_windex & 6'h3a == pht_waddr ? pht_2_58 : _GEN_2873; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2875 = 3'h2 == pht_windex & 6'h3b == pht_waddr ? pht_2_59 : _GEN_2874; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2876 = 3'h2 == pht_windex & 6'h3c == pht_waddr ? pht_2_60 : _GEN_2875; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2877 = 3'h2 == pht_windex & 6'h3d == pht_waddr ? pht_2_61 : _GEN_2876; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2878 = 3'h2 == pht_windex & 6'h3e == pht_waddr ? pht_2_62 : _GEN_2877; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2879 = 3'h2 == pht_windex & 6'h3f == pht_waddr ? pht_2_63 : _GEN_2878; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2880 = 3'h2 == pht_windex & 7'h40 == _GEN_14784 ? pht_2_64 : _GEN_2879; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2881 = 3'h2 == pht_windex & 7'h41 == _GEN_14784 ? pht_2_65 : _GEN_2880; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2882 = 3'h2 == pht_windex & 7'h42 == _GEN_14784 ? pht_2_66 : _GEN_2881; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2883 = 3'h2 == pht_windex & 7'h43 == _GEN_14784 ? pht_2_67 : _GEN_2882; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2884 = 3'h2 == pht_windex & 7'h44 == _GEN_14784 ? pht_2_68 : _GEN_2883; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2885 = 3'h2 == pht_windex & 7'h45 == _GEN_14784 ? pht_2_69 : _GEN_2884; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2886 = 3'h2 == pht_windex & 7'h46 == _GEN_14784 ? pht_2_70 : _GEN_2885; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2887 = 3'h2 == pht_windex & 7'h47 == _GEN_14784 ? pht_2_71 : _GEN_2886; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2888 = 3'h2 == pht_windex & 7'h48 == _GEN_14784 ? pht_2_72 : _GEN_2887; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2889 = 3'h2 == pht_windex & 7'h49 == _GEN_14784 ? pht_2_73 : _GEN_2888; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2890 = 3'h2 == pht_windex & 7'h4a == _GEN_14784 ? pht_2_74 : _GEN_2889; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2891 = 3'h2 == pht_windex & 7'h4b == _GEN_14784 ? pht_2_75 : _GEN_2890; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2892 = 3'h2 == pht_windex & 7'h4c == _GEN_14784 ? pht_2_76 : _GEN_2891; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2893 = 3'h2 == pht_windex & 7'h4d == _GEN_14784 ? pht_2_77 : _GEN_2892; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2894 = 3'h2 == pht_windex & 7'h4e == _GEN_14784 ? pht_2_78 : _GEN_2893; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2895 = 3'h2 == pht_windex & 7'h4f == _GEN_14784 ? pht_2_79 : _GEN_2894; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2896 = 3'h2 == pht_windex & 7'h50 == _GEN_14784 ? pht_2_80 : _GEN_2895; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2897 = 3'h2 == pht_windex & 7'h51 == _GEN_14784 ? pht_2_81 : _GEN_2896; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2898 = 3'h2 == pht_windex & 7'h52 == _GEN_14784 ? pht_2_82 : _GEN_2897; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2899 = 3'h2 == pht_windex & 7'h53 == _GEN_14784 ? pht_2_83 : _GEN_2898; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2900 = 3'h2 == pht_windex & 7'h54 == _GEN_14784 ? pht_2_84 : _GEN_2899; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2901 = 3'h2 == pht_windex & 7'h55 == _GEN_14784 ? pht_2_85 : _GEN_2900; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2902 = 3'h2 == pht_windex & 7'h56 == _GEN_14784 ? pht_2_86 : _GEN_2901; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2903 = 3'h2 == pht_windex & 7'h57 == _GEN_14784 ? pht_2_87 : _GEN_2902; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2904 = 3'h2 == pht_windex & 7'h58 == _GEN_14784 ? pht_2_88 : _GEN_2903; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2905 = 3'h2 == pht_windex & 7'h59 == _GEN_14784 ? pht_2_89 : _GEN_2904; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2906 = 3'h2 == pht_windex & 7'h5a == _GEN_14784 ? pht_2_90 : _GEN_2905; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2907 = 3'h2 == pht_windex & 7'h5b == _GEN_14784 ? pht_2_91 : _GEN_2906; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2908 = 3'h2 == pht_windex & 7'h5c == _GEN_14784 ? pht_2_92 : _GEN_2907; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2909 = 3'h2 == pht_windex & 7'h5d == _GEN_14784 ? pht_2_93 : _GEN_2908; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2910 = 3'h2 == pht_windex & 7'h5e == _GEN_14784 ? pht_2_94 : _GEN_2909; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2911 = 3'h2 == pht_windex & 7'h5f == _GEN_14784 ? pht_2_95 : _GEN_2910; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2912 = 3'h2 == pht_windex & 7'h60 == _GEN_14784 ? pht_2_96 : _GEN_2911; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2913 = 3'h2 == pht_windex & 7'h61 == _GEN_14784 ? pht_2_97 : _GEN_2912; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2914 = 3'h2 == pht_windex & 7'h62 == _GEN_14784 ? pht_2_98 : _GEN_2913; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2915 = 3'h2 == pht_windex & 7'h63 == _GEN_14784 ? pht_2_99 : _GEN_2914; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2916 = 3'h2 == pht_windex & 7'h64 == _GEN_14784 ? pht_2_100 : _GEN_2915; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2917 = 3'h2 == pht_windex & 7'h65 == _GEN_14784 ? pht_2_101 : _GEN_2916; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2918 = 3'h2 == pht_windex & 7'h66 == _GEN_14784 ? pht_2_102 : _GEN_2917; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2919 = 3'h2 == pht_windex & 7'h67 == _GEN_14784 ? pht_2_103 : _GEN_2918; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2920 = 3'h2 == pht_windex & 7'h68 == _GEN_14784 ? pht_2_104 : _GEN_2919; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2921 = 3'h2 == pht_windex & 7'h69 == _GEN_14784 ? pht_2_105 : _GEN_2920; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2922 = 3'h2 == pht_windex & 7'h6a == _GEN_14784 ? pht_2_106 : _GEN_2921; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2923 = 3'h2 == pht_windex & 7'h6b == _GEN_14784 ? pht_2_107 : _GEN_2922; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2924 = 3'h2 == pht_windex & 7'h6c == _GEN_14784 ? pht_2_108 : _GEN_2923; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2925 = 3'h2 == pht_windex & 7'h6d == _GEN_14784 ? pht_2_109 : _GEN_2924; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2926 = 3'h2 == pht_windex & 7'h6e == _GEN_14784 ? pht_2_110 : _GEN_2925; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2927 = 3'h2 == pht_windex & 7'h6f == _GEN_14784 ? pht_2_111 : _GEN_2926; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2928 = 3'h2 == pht_windex & 7'h70 == _GEN_14784 ? pht_2_112 : _GEN_2927; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2929 = 3'h2 == pht_windex & 7'h71 == _GEN_14784 ? pht_2_113 : _GEN_2928; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2930 = 3'h2 == pht_windex & 7'h72 == _GEN_14784 ? pht_2_114 : _GEN_2929; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2931 = 3'h2 == pht_windex & 7'h73 == _GEN_14784 ? pht_2_115 : _GEN_2930; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2932 = 3'h2 == pht_windex & 7'h74 == _GEN_14784 ? pht_2_116 : _GEN_2931; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2933 = 3'h2 == pht_windex & 7'h75 == _GEN_14784 ? pht_2_117 : _GEN_2932; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2934 = 3'h2 == pht_windex & 7'h76 == _GEN_14784 ? pht_2_118 : _GEN_2933; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2935 = 3'h2 == pht_windex & 7'h77 == _GEN_14784 ? pht_2_119 : _GEN_2934; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2936 = 3'h2 == pht_windex & 7'h78 == _GEN_14784 ? pht_2_120 : _GEN_2935; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2937 = 3'h2 == pht_windex & 7'h79 == _GEN_14784 ? pht_2_121 : _GEN_2936; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2938 = 3'h2 == pht_windex & 7'h7a == _GEN_14784 ? pht_2_122 : _GEN_2937; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2939 = 3'h2 == pht_windex & 7'h7b == _GEN_14784 ? pht_2_123 : _GEN_2938; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2940 = 3'h2 == pht_windex & 7'h7c == _GEN_14784 ? pht_2_124 : _GEN_2939; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2941 = 3'h2 == pht_windex & 7'h7d == _GEN_14784 ? pht_2_125 : _GEN_2940; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2942 = 3'h2 == pht_windex & 7'h7e == _GEN_14784 ? pht_2_126 : _GEN_2941; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2943 = 3'h2 == pht_windex & 7'h7f == _GEN_14784 ? pht_2_127 : _GEN_2942; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2944 = 3'h2 == pht_windex & 8'h80 == _GEN_14976 ? pht_2_128 : _GEN_2943; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2945 = 3'h2 == pht_windex & 8'h81 == _GEN_14976 ? pht_2_129 : _GEN_2944; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2946 = 3'h2 == pht_windex & 8'h82 == _GEN_14976 ? pht_2_130 : _GEN_2945; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2947 = 3'h2 == pht_windex & 8'h83 == _GEN_14976 ? pht_2_131 : _GEN_2946; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2948 = 3'h2 == pht_windex & 8'h84 == _GEN_14976 ? pht_2_132 : _GEN_2947; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2949 = 3'h2 == pht_windex & 8'h85 == _GEN_14976 ? pht_2_133 : _GEN_2948; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2950 = 3'h2 == pht_windex & 8'h86 == _GEN_14976 ? pht_2_134 : _GEN_2949; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2951 = 3'h2 == pht_windex & 8'h87 == _GEN_14976 ? pht_2_135 : _GEN_2950; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2952 = 3'h2 == pht_windex & 8'h88 == _GEN_14976 ? pht_2_136 : _GEN_2951; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2953 = 3'h2 == pht_windex & 8'h89 == _GEN_14976 ? pht_2_137 : _GEN_2952; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2954 = 3'h2 == pht_windex & 8'h8a == _GEN_14976 ? pht_2_138 : _GEN_2953; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2955 = 3'h2 == pht_windex & 8'h8b == _GEN_14976 ? pht_2_139 : _GEN_2954; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2956 = 3'h2 == pht_windex & 8'h8c == _GEN_14976 ? pht_2_140 : _GEN_2955; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2957 = 3'h2 == pht_windex & 8'h8d == _GEN_14976 ? pht_2_141 : _GEN_2956; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2958 = 3'h2 == pht_windex & 8'h8e == _GEN_14976 ? pht_2_142 : _GEN_2957; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2959 = 3'h2 == pht_windex & 8'h8f == _GEN_14976 ? pht_2_143 : _GEN_2958; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2960 = 3'h2 == pht_windex & 8'h90 == _GEN_14976 ? pht_2_144 : _GEN_2959; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2961 = 3'h2 == pht_windex & 8'h91 == _GEN_14976 ? pht_2_145 : _GEN_2960; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2962 = 3'h2 == pht_windex & 8'h92 == _GEN_14976 ? pht_2_146 : _GEN_2961; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2963 = 3'h2 == pht_windex & 8'h93 == _GEN_14976 ? pht_2_147 : _GEN_2962; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2964 = 3'h2 == pht_windex & 8'h94 == _GEN_14976 ? pht_2_148 : _GEN_2963; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2965 = 3'h2 == pht_windex & 8'h95 == _GEN_14976 ? pht_2_149 : _GEN_2964; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2966 = 3'h2 == pht_windex & 8'h96 == _GEN_14976 ? pht_2_150 : _GEN_2965; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2967 = 3'h2 == pht_windex & 8'h97 == _GEN_14976 ? pht_2_151 : _GEN_2966; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2968 = 3'h2 == pht_windex & 8'h98 == _GEN_14976 ? pht_2_152 : _GEN_2967; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2969 = 3'h2 == pht_windex & 8'h99 == _GEN_14976 ? pht_2_153 : _GEN_2968; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2970 = 3'h2 == pht_windex & 8'h9a == _GEN_14976 ? pht_2_154 : _GEN_2969; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2971 = 3'h2 == pht_windex & 8'h9b == _GEN_14976 ? pht_2_155 : _GEN_2970; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2972 = 3'h2 == pht_windex & 8'h9c == _GEN_14976 ? pht_2_156 : _GEN_2971; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2973 = 3'h2 == pht_windex & 8'h9d == _GEN_14976 ? pht_2_157 : _GEN_2972; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2974 = 3'h2 == pht_windex & 8'h9e == _GEN_14976 ? pht_2_158 : _GEN_2973; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2975 = 3'h2 == pht_windex & 8'h9f == _GEN_14976 ? pht_2_159 : _GEN_2974; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2976 = 3'h2 == pht_windex & 8'ha0 == _GEN_14976 ? pht_2_160 : _GEN_2975; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2977 = 3'h2 == pht_windex & 8'ha1 == _GEN_14976 ? pht_2_161 : _GEN_2976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2978 = 3'h2 == pht_windex & 8'ha2 == _GEN_14976 ? pht_2_162 : _GEN_2977; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2979 = 3'h2 == pht_windex & 8'ha3 == _GEN_14976 ? pht_2_163 : _GEN_2978; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2980 = 3'h2 == pht_windex & 8'ha4 == _GEN_14976 ? pht_2_164 : _GEN_2979; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2981 = 3'h2 == pht_windex & 8'ha5 == _GEN_14976 ? pht_2_165 : _GEN_2980; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2982 = 3'h2 == pht_windex & 8'ha6 == _GEN_14976 ? pht_2_166 : _GEN_2981; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2983 = 3'h2 == pht_windex & 8'ha7 == _GEN_14976 ? pht_2_167 : _GEN_2982; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2984 = 3'h2 == pht_windex & 8'ha8 == _GEN_14976 ? pht_2_168 : _GEN_2983; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2985 = 3'h2 == pht_windex & 8'ha9 == _GEN_14976 ? pht_2_169 : _GEN_2984; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2986 = 3'h2 == pht_windex & 8'haa == _GEN_14976 ? pht_2_170 : _GEN_2985; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2987 = 3'h2 == pht_windex & 8'hab == _GEN_14976 ? pht_2_171 : _GEN_2986; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2988 = 3'h2 == pht_windex & 8'hac == _GEN_14976 ? pht_2_172 : _GEN_2987; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2989 = 3'h2 == pht_windex & 8'had == _GEN_14976 ? pht_2_173 : _GEN_2988; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2990 = 3'h2 == pht_windex & 8'hae == _GEN_14976 ? pht_2_174 : _GEN_2989; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2991 = 3'h2 == pht_windex & 8'haf == _GEN_14976 ? pht_2_175 : _GEN_2990; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2992 = 3'h2 == pht_windex & 8'hb0 == _GEN_14976 ? pht_2_176 : _GEN_2991; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2993 = 3'h2 == pht_windex & 8'hb1 == _GEN_14976 ? pht_2_177 : _GEN_2992; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2994 = 3'h2 == pht_windex & 8'hb2 == _GEN_14976 ? pht_2_178 : _GEN_2993; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2995 = 3'h2 == pht_windex & 8'hb3 == _GEN_14976 ? pht_2_179 : _GEN_2994; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2996 = 3'h2 == pht_windex & 8'hb4 == _GEN_14976 ? pht_2_180 : _GEN_2995; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2997 = 3'h2 == pht_windex & 8'hb5 == _GEN_14976 ? pht_2_181 : _GEN_2996; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2998 = 3'h2 == pht_windex & 8'hb6 == _GEN_14976 ? pht_2_182 : _GEN_2997; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_2999 = 3'h2 == pht_windex & 8'hb7 == _GEN_14976 ? pht_2_183 : _GEN_2998; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3000 = 3'h2 == pht_windex & 8'hb8 == _GEN_14976 ? pht_2_184 : _GEN_2999; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3001 = 3'h2 == pht_windex & 8'hb9 == _GEN_14976 ? pht_2_185 : _GEN_3000; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3002 = 3'h2 == pht_windex & 8'hba == _GEN_14976 ? pht_2_186 : _GEN_3001; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3003 = 3'h2 == pht_windex & 8'hbb == _GEN_14976 ? pht_2_187 : _GEN_3002; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3004 = 3'h2 == pht_windex & 8'hbc == _GEN_14976 ? pht_2_188 : _GEN_3003; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3005 = 3'h2 == pht_windex & 8'hbd == _GEN_14976 ? pht_2_189 : _GEN_3004; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3006 = 3'h2 == pht_windex & 8'hbe == _GEN_14976 ? pht_2_190 : _GEN_3005; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3007 = 3'h2 == pht_windex & 8'hbf == _GEN_14976 ? pht_2_191 : _GEN_3006; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3008 = 3'h2 == pht_windex & 8'hc0 == _GEN_14976 ? pht_2_192 : _GEN_3007; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3009 = 3'h2 == pht_windex & 8'hc1 == _GEN_14976 ? pht_2_193 : _GEN_3008; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3010 = 3'h2 == pht_windex & 8'hc2 == _GEN_14976 ? pht_2_194 : _GEN_3009; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3011 = 3'h2 == pht_windex & 8'hc3 == _GEN_14976 ? pht_2_195 : _GEN_3010; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3012 = 3'h2 == pht_windex & 8'hc4 == _GEN_14976 ? pht_2_196 : _GEN_3011; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3013 = 3'h2 == pht_windex & 8'hc5 == _GEN_14976 ? pht_2_197 : _GEN_3012; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3014 = 3'h2 == pht_windex & 8'hc6 == _GEN_14976 ? pht_2_198 : _GEN_3013; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3015 = 3'h2 == pht_windex & 8'hc7 == _GEN_14976 ? pht_2_199 : _GEN_3014; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3016 = 3'h2 == pht_windex & 8'hc8 == _GEN_14976 ? pht_2_200 : _GEN_3015; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3017 = 3'h2 == pht_windex & 8'hc9 == _GEN_14976 ? pht_2_201 : _GEN_3016; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3018 = 3'h2 == pht_windex & 8'hca == _GEN_14976 ? pht_2_202 : _GEN_3017; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3019 = 3'h2 == pht_windex & 8'hcb == _GEN_14976 ? pht_2_203 : _GEN_3018; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3020 = 3'h2 == pht_windex & 8'hcc == _GEN_14976 ? pht_2_204 : _GEN_3019; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3021 = 3'h2 == pht_windex & 8'hcd == _GEN_14976 ? pht_2_205 : _GEN_3020; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3022 = 3'h2 == pht_windex & 8'hce == _GEN_14976 ? pht_2_206 : _GEN_3021; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3023 = 3'h2 == pht_windex & 8'hcf == _GEN_14976 ? pht_2_207 : _GEN_3022; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3024 = 3'h2 == pht_windex & 8'hd0 == _GEN_14976 ? pht_2_208 : _GEN_3023; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3025 = 3'h2 == pht_windex & 8'hd1 == _GEN_14976 ? pht_2_209 : _GEN_3024; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3026 = 3'h2 == pht_windex & 8'hd2 == _GEN_14976 ? pht_2_210 : _GEN_3025; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3027 = 3'h2 == pht_windex & 8'hd3 == _GEN_14976 ? pht_2_211 : _GEN_3026; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3028 = 3'h2 == pht_windex & 8'hd4 == _GEN_14976 ? pht_2_212 : _GEN_3027; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3029 = 3'h2 == pht_windex & 8'hd5 == _GEN_14976 ? pht_2_213 : _GEN_3028; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3030 = 3'h2 == pht_windex & 8'hd6 == _GEN_14976 ? pht_2_214 : _GEN_3029; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3031 = 3'h2 == pht_windex & 8'hd7 == _GEN_14976 ? pht_2_215 : _GEN_3030; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3032 = 3'h2 == pht_windex & 8'hd8 == _GEN_14976 ? pht_2_216 : _GEN_3031; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3033 = 3'h2 == pht_windex & 8'hd9 == _GEN_14976 ? pht_2_217 : _GEN_3032; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3034 = 3'h2 == pht_windex & 8'hda == _GEN_14976 ? pht_2_218 : _GEN_3033; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3035 = 3'h2 == pht_windex & 8'hdb == _GEN_14976 ? pht_2_219 : _GEN_3034; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3036 = 3'h2 == pht_windex & 8'hdc == _GEN_14976 ? pht_2_220 : _GEN_3035; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3037 = 3'h2 == pht_windex & 8'hdd == _GEN_14976 ? pht_2_221 : _GEN_3036; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3038 = 3'h2 == pht_windex & 8'hde == _GEN_14976 ? pht_2_222 : _GEN_3037; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3039 = 3'h2 == pht_windex & 8'hdf == _GEN_14976 ? pht_2_223 : _GEN_3038; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3040 = 3'h2 == pht_windex & 8'he0 == _GEN_14976 ? pht_2_224 : _GEN_3039; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3041 = 3'h2 == pht_windex & 8'he1 == _GEN_14976 ? pht_2_225 : _GEN_3040; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3042 = 3'h2 == pht_windex & 8'he2 == _GEN_14976 ? pht_2_226 : _GEN_3041; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3043 = 3'h2 == pht_windex & 8'he3 == _GEN_14976 ? pht_2_227 : _GEN_3042; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3044 = 3'h2 == pht_windex & 8'he4 == _GEN_14976 ? pht_2_228 : _GEN_3043; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3045 = 3'h2 == pht_windex & 8'he5 == _GEN_14976 ? pht_2_229 : _GEN_3044; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3046 = 3'h2 == pht_windex & 8'he6 == _GEN_14976 ? pht_2_230 : _GEN_3045; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3047 = 3'h2 == pht_windex & 8'he7 == _GEN_14976 ? pht_2_231 : _GEN_3046; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3048 = 3'h2 == pht_windex & 8'he8 == _GEN_14976 ? pht_2_232 : _GEN_3047; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3049 = 3'h2 == pht_windex & 8'he9 == _GEN_14976 ? pht_2_233 : _GEN_3048; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3050 = 3'h2 == pht_windex & 8'hea == _GEN_14976 ? pht_2_234 : _GEN_3049; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3051 = 3'h2 == pht_windex & 8'heb == _GEN_14976 ? pht_2_235 : _GEN_3050; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3052 = 3'h2 == pht_windex & 8'hec == _GEN_14976 ? pht_2_236 : _GEN_3051; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3053 = 3'h2 == pht_windex & 8'hed == _GEN_14976 ? pht_2_237 : _GEN_3052; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3054 = 3'h2 == pht_windex & 8'hee == _GEN_14976 ? pht_2_238 : _GEN_3053; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3055 = 3'h2 == pht_windex & 8'hef == _GEN_14976 ? pht_2_239 : _GEN_3054; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3056 = 3'h2 == pht_windex & 8'hf0 == _GEN_14976 ? pht_2_240 : _GEN_3055; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3057 = 3'h2 == pht_windex & 8'hf1 == _GEN_14976 ? pht_2_241 : _GEN_3056; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3058 = 3'h2 == pht_windex & 8'hf2 == _GEN_14976 ? pht_2_242 : _GEN_3057; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3059 = 3'h2 == pht_windex & 8'hf3 == _GEN_14976 ? pht_2_243 : _GEN_3058; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3060 = 3'h2 == pht_windex & 8'hf4 == _GEN_14976 ? pht_2_244 : _GEN_3059; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3061 = 3'h2 == pht_windex & 8'hf5 == _GEN_14976 ? pht_2_245 : _GEN_3060; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3062 = 3'h2 == pht_windex & 8'hf6 == _GEN_14976 ? pht_2_246 : _GEN_3061; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3063 = 3'h2 == pht_windex & 8'hf7 == _GEN_14976 ? pht_2_247 : _GEN_3062; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3064 = 3'h2 == pht_windex & 8'hf8 == _GEN_14976 ? pht_2_248 : _GEN_3063; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3065 = 3'h2 == pht_windex & 8'hf9 == _GEN_14976 ? pht_2_249 : _GEN_3064; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3066 = 3'h2 == pht_windex & 8'hfa == _GEN_14976 ? pht_2_250 : _GEN_3065; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3067 = 3'h2 == pht_windex & 8'hfb == _GEN_14976 ? pht_2_251 : _GEN_3066; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3068 = 3'h2 == pht_windex & 8'hfc == _GEN_14976 ? pht_2_252 : _GEN_3067; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3069 = 3'h2 == pht_windex & 8'hfd == _GEN_14976 ? pht_2_253 : _GEN_3068; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3070 = 3'h2 == pht_windex & 8'hfe == _GEN_14976 ? pht_2_254 : _GEN_3069; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3071 = 3'h2 == pht_windex & 8'hff == _GEN_14976 ? pht_2_255 : _GEN_3070; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_16768 = 3'h3 == pht_windex; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3072 = 3'h3 == pht_windex & 6'h0 == pht_waddr ? pht_3_0 : _GEN_3071; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3073 = 3'h3 == pht_windex & 6'h1 == pht_waddr ? pht_3_1 : _GEN_3072; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3074 = 3'h3 == pht_windex & 6'h2 == pht_waddr ? pht_3_2 : _GEN_3073; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3075 = 3'h3 == pht_windex & 6'h3 == pht_waddr ? pht_3_3 : _GEN_3074; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3076 = 3'h3 == pht_windex & 6'h4 == pht_waddr ? pht_3_4 : _GEN_3075; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3077 = 3'h3 == pht_windex & 6'h5 == pht_waddr ? pht_3_5 : _GEN_3076; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3078 = 3'h3 == pht_windex & 6'h6 == pht_waddr ? pht_3_6 : _GEN_3077; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3079 = 3'h3 == pht_windex & 6'h7 == pht_waddr ? pht_3_7 : _GEN_3078; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3080 = 3'h3 == pht_windex & 6'h8 == pht_waddr ? pht_3_8 : _GEN_3079; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3081 = 3'h3 == pht_windex & 6'h9 == pht_waddr ? pht_3_9 : _GEN_3080; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3082 = 3'h3 == pht_windex & 6'ha == pht_waddr ? pht_3_10 : _GEN_3081; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3083 = 3'h3 == pht_windex & 6'hb == pht_waddr ? pht_3_11 : _GEN_3082; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3084 = 3'h3 == pht_windex & 6'hc == pht_waddr ? pht_3_12 : _GEN_3083; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3085 = 3'h3 == pht_windex & 6'hd == pht_waddr ? pht_3_13 : _GEN_3084; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3086 = 3'h3 == pht_windex & 6'he == pht_waddr ? pht_3_14 : _GEN_3085; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3087 = 3'h3 == pht_windex & 6'hf == pht_waddr ? pht_3_15 : _GEN_3086; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3088 = 3'h3 == pht_windex & 6'h10 == pht_waddr ? pht_3_16 : _GEN_3087; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3089 = 3'h3 == pht_windex & 6'h11 == pht_waddr ? pht_3_17 : _GEN_3088; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3090 = 3'h3 == pht_windex & 6'h12 == pht_waddr ? pht_3_18 : _GEN_3089; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3091 = 3'h3 == pht_windex & 6'h13 == pht_waddr ? pht_3_19 : _GEN_3090; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3092 = 3'h3 == pht_windex & 6'h14 == pht_waddr ? pht_3_20 : _GEN_3091; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3093 = 3'h3 == pht_windex & 6'h15 == pht_waddr ? pht_3_21 : _GEN_3092; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3094 = 3'h3 == pht_windex & 6'h16 == pht_waddr ? pht_3_22 : _GEN_3093; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3095 = 3'h3 == pht_windex & 6'h17 == pht_waddr ? pht_3_23 : _GEN_3094; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3096 = 3'h3 == pht_windex & 6'h18 == pht_waddr ? pht_3_24 : _GEN_3095; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3097 = 3'h3 == pht_windex & 6'h19 == pht_waddr ? pht_3_25 : _GEN_3096; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3098 = 3'h3 == pht_windex & 6'h1a == pht_waddr ? pht_3_26 : _GEN_3097; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3099 = 3'h3 == pht_windex & 6'h1b == pht_waddr ? pht_3_27 : _GEN_3098; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3100 = 3'h3 == pht_windex & 6'h1c == pht_waddr ? pht_3_28 : _GEN_3099; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3101 = 3'h3 == pht_windex & 6'h1d == pht_waddr ? pht_3_29 : _GEN_3100; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3102 = 3'h3 == pht_windex & 6'h1e == pht_waddr ? pht_3_30 : _GEN_3101; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3103 = 3'h3 == pht_windex & 6'h1f == pht_waddr ? pht_3_31 : _GEN_3102; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3104 = 3'h3 == pht_windex & 6'h20 == pht_waddr ? pht_3_32 : _GEN_3103; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3105 = 3'h3 == pht_windex & 6'h21 == pht_waddr ? pht_3_33 : _GEN_3104; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3106 = 3'h3 == pht_windex & 6'h22 == pht_waddr ? pht_3_34 : _GEN_3105; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3107 = 3'h3 == pht_windex & 6'h23 == pht_waddr ? pht_3_35 : _GEN_3106; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3108 = 3'h3 == pht_windex & 6'h24 == pht_waddr ? pht_3_36 : _GEN_3107; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3109 = 3'h3 == pht_windex & 6'h25 == pht_waddr ? pht_3_37 : _GEN_3108; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3110 = 3'h3 == pht_windex & 6'h26 == pht_waddr ? pht_3_38 : _GEN_3109; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3111 = 3'h3 == pht_windex & 6'h27 == pht_waddr ? pht_3_39 : _GEN_3110; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3112 = 3'h3 == pht_windex & 6'h28 == pht_waddr ? pht_3_40 : _GEN_3111; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3113 = 3'h3 == pht_windex & 6'h29 == pht_waddr ? pht_3_41 : _GEN_3112; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3114 = 3'h3 == pht_windex & 6'h2a == pht_waddr ? pht_3_42 : _GEN_3113; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3115 = 3'h3 == pht_windex & 6'h2b == pht_waddr ? pht_3_43 : _GEN_3114; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3116 = 3'h3 == pht_windex & 6'h2c == pht_waddr ? pht_3_44 : _GEN_3115; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3117 = 3'h3 == pht_windex & 6'h2d == pht_waddr ? pht_3_45 : _GEN_3116; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3118 = 3'h3 == pht_windex & 6'h2e == pht_waddr ? pht_3_46 : _GEN_3117; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3119 = 3'h3 == pht_windex & 6'h2f == pht_waddr ? pht_3_47 : _GEN_3118; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3120 = 3'h3 == pht_windex & 6'h30 == pht_waddr ? pht_3_48 : _GEN_3119; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3121 = 3'h3 == pht_windex & 6'h31 == pht_waddr ? pht_3_49 : _GEN_3120; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3122 = 3'h3 == pht_windex & 6'h32 == pht_waddr ? pht_3_50 : _GEN_3121; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3123 = 3'h3 == pht_windex & 6'h33 == pht_waddr ? pht_3_51 : _GEN_3122; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3124 = 3'h3 == pht_windex & 6'h34 == pht_waddr ? pht_3_52 : _GEN_3123; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3125 = 3'h3 == pht_windex & 6'h35 == pht_waddr ? pht_3_53 : _GEN_3124; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3126 = 3'h3 == pht_windex & 6'h36 == pht_waddr ? pht_3_54 : _GEN_3125; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3127 = 3'h3 == pht_windex & 6'h37 == pht_waddr ? pht_3_55 : _GEN_3126; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3128 = 3'h3 == pht_windex & 6'h38 == pht_waddr ? pht_3_56 : _GEN_3127; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3129 = 3'h3 == pht_windex & 6'h39 == pht_waddr ? pht_3_57 : _GEN_3128; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3130 = 3'h3 == pht_windex & 6'h3a == pht_waddr ? pht_3_58 : _GEN_3129; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3131 = 3'h3 == pht_windex & 6'h3b == pht_waddr ? pht_3_59 : _GEN_3130; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3132 = 3'h3 == pht_windex & 6'h3c == pht_waddr ? pht_3_60 : _GEN_3131; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3133 = 3'h3 == pht_windex & 6'h3d == pht_waddr ? pht_3_61 : _GEN_3132; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3134 = 3'h3 == pht_windex & 6'h3e == pht_waddr ? pht_3_62 : _GEN_3133; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3135 = 3'h3 == pht_windex & 6'h3f == pht_waddr ? pht_3_63 : _GEN_3134; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3136 = 3'h3 == pht_windex & 7'h40 == _GEN_14784 ? pht_3_64 : _GEN_3135; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3137 = 3'h3 == pht_windex & 7'h41 == _GEN_14784 ? pht_3_65 : _GEN_3136; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3138 = 3'h3 == pht_windex & 7'h42 == _GEN_14784 ? pht_3_66 : _GEN_3137; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3139 = 3'h3 == pht_windex & 7'h43 == _GEN_14784 ? pht_3_67 : _GEN_3138; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3140 = 3'h3 == pht_windex & 7'h44 == _GEN_14784 ? pht_3_68 : _GEN_3139; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3141 = 3'h3 == pht_windex & 7'h45 == _GEN_14784 ? pht_3_69 : _GEN_3140; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3142 = 3'h3 == pht_windex & 7'h46 == _GEN_14784 ? pht_3_70 : _GEN_3141; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3143 = 3'h3 == pht_windex & 7'h47 == _GEN_14784 ? pht_3_71 : _GEN_3142; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3144 = 3'h3 == pht_windex & 7'h48 == _GEN_14784 ? pht_3_72 : _GEN_3143; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3145 = 3'h3 == pht_windex & 7'h49 == _GEN_14784 ? pht_3_73 : _GEN_3144; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3146 = 3'h3 == pht_windex & 7'h4a == _GEN_14784 ? pht_3_74 : _GEN_3145; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3147 = 3'h3 == pht_windex & 7'h4b == _GEN_14784 ? pht_3_75 : _GEN_3146; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3148 = 3'h3 == pht_windex & 7'h4c == _GEN_14784 ? pht_3_76 : _GEN_3147; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3149 = 3'h3 == pht_windex & 7'h4d == _GEN_14784 ? pht_3_77 : _GEN_3148; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3150 = 3'h3 == pht_windex & 7'h4e == _GEN_14784 ? pht_3_78 : _GEN_3149; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3151 = 3'h3 == pht_windex & 7'h4f == _GEN_14784 ? pht_3_79 : _GEN_3150; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3152 = 3'h3 == pht_windex & 7'h50 == _GEN_14784 ? pht_3_80 : _GEN_3151; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3153 = 3'h3 == pht_windex & 7'h51 == _GEN_14784 ? pht_3_81 : _GEN_3152; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3154 = 3'h3 == pht_windex & 7'h52 == _GEN_14784 ? pht_3_82 : _GEN_3153; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3155 = 3'h3 == pht_windex & 7'h53 == _GEN_14784 ? pht_3_83 : _GEN_3154; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3156 = 3'h3 == pht_windex & 7'h54 == _GEN_14784 ? pht_3_84 : _GEN_3155; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3157 = 3'h3 == pht_windex & 7'h55 == _GEN_14784 ? pht_3_85 : _GEN_3156; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3158 = 3'h3 == pht_windex & 7'h56 == _GEN_14784 ? pht_3_86 : _GEN_3157; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3159 = 3'h3 == pht_windex & 7'h57 == _GEN_14784 ? pht_3_87 : _GEN_3158; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3160 = 3'h3 == pht_windex & 7'h58 == _GEN_14784 ? pht_3_88 : _GEN_3159; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3161 = 3'h3 == pht_windex & 7'h59 == _GEN_14784 ? pht_3_89 : _GEN_3160; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3162 = 3'h3 == pht_windex & 7'h5a == _GEN_14784 ? pht_3_90 : _GEN_3161; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3163 = 3'h3 == pht_windex & 7'h5b == _GEN_14784 ? pht_3_91 : _GEN_3162; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3164 = 3'h3 == pht_windex & 7'h5c == _GEN_14784 ? pht_3_92 : _GEN_3163; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3165 = 3'h3 == pht_windex & 7'h5d == _GEN_14784 ? pht_3_93 : _GEN_3164; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3166 = 3'h3 == pht_windex & 7'h5e == _GEN_14784 ? pht_3_94 : _GEN_3165; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3167 = 3'h3 == pht_windex & 7'h5f == _GEN_14784 ? pht_3_95 : _GEN_3166; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3168 = 3'h3 == pht_windex & 7'h60 == _GEN_14784 ? pht_3_96 : _GEN_3167; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3169 = 3'h3 == pht_windex & 7'h61 == _GEN_14784 ? pht_3_97 : _GEN_3168; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3170 = 3'h3 == pht_windex & 7'h62 == _GEN_14784 ? pht_3_98 : _GEN_3169; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3171 = 3'h3 == pht_windex & 7'h63 == _GEN_14784 ? pht_3_99 : _GEN_3170; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3172 = 3'h3 == pht_windex & 7'h64 == _GEN_14784 ? pht_3_100 : _GEN_3171; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3173 = 3'h3 == pht_windex & 7'h65 == _GEN_14784 ? pht_3_101 : _GEN_3172; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3174 = 3'h3 == pht_windex & 7'h66 == _GEN_14784 ? pht_3_102 : _GEN_3173; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3175 = 3'h3 == pht_windex & 7'h67 == _GEN_14784 ? pht_3_103 : _GEN_3174; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3176 = 3'h3 == pht_windex & 7'h68 == _GEN_14784 ? pht_3_104 : _GEN_3175; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3177 = 3'h3 == pht_windex & 7'h69 == _GEN_14784 ? pht_3_105 : _GEN_3176; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3178 = 3'h3 == pht_windex & 7'h6a == _GEN_14784 ? pht_3_106 : _GEN_3177; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3179 = 3'h3 == pht_windex & 7'h6b == _GEN_14784 ? pht_3_107 : _GEN_3178; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3180 = 3'h3 == pht_windex & 7'h6c == _GEN_14784 ? pht_3_108 : _GEN_3179; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3181 = 3'h3 == pht_windex & 7'h6d == _GEN_14784 ? pht_3_109 : _GEN_3180; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3182 = 3'h3 == pht_windex & 7'h6e == _GEN_14784 ? pht_3_110 : _GEN_3181; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3183 = 3'h3 == pht_windex & 7'h6f == _GEN_14784 ? pht_3_111 : _GEN_3182; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3184 = 3'h3 == pht_windex & 7'h70 == _GEN_14784 ? pht_3_112 : _GEN_3183; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3185 = 3'h3 == pht_windex & 7'h71 == _GEN_14784 ? pht_3_113 : _GEN_3184; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3186 = 3'h3 == pht_windex & 7'h72 == _GEN_14784 ? pht_3_114 : _GEN_3185; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3187 = 3'h3 == pht_windex & 7'h73 == _GEN_14784 ? pht_3_115 : _GEN_3186; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3188 = 3'h3 == pht_windex & 7'h74 == _GEN_14784 ? pht_3_116 : _GEN_3187; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3189 = 3'h3 == pht_windex & 7'h75 == _GEN_14784 ? pht_3_117 : _GEN_3188; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3190 = 3'h3 == pht_windex & 7'h76 == _GEN_14784 ? pht_3_118 : _GEN_3189; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3191 = 3'h3 == pht_windex & 7'h77 == _GEN_14784 ? pht_3_119 : _GEN_3190; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3192 = 3'h3 == pht_windex & 7'h78 == _GEN_14784 ? pht_3_120 : _GEN_3191; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3193 = 3'h3 == pht_windex & 7'h79 == _GEN_14784 ? pht_3_121 : _GEN_3192; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3194 = 3'h3 == pht_windex & 7'h7a == _GEN_14784 ? pht_3_122 : _GEN_3193; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3195 = 3'h3 == pht_windex & 7'h7b == _GEN_14784 ? pht_3_123 : _GEN_3194; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3196 = 3'h3 == pht_windex & 7'h7c == _GEN_14784 ? pht_3_124 : _GEN_3195; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3197 = 3'h3 == pht_windex & 7'h7d == _GEN_14784 ? pht_3_125 : _GEN_3196; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3198 = 3'h3 == pht_windex & 7'h7e == _GEN_14784 ? pht_3_126 : _GEN_3197; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3199 = 3'h3 == pht_windex & 7'h7f == _GEN_14784 ? pht_3_127 : _GEN_3198; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3200 = 3'h3 == pht_windex & 8'h80 == _GEN_14976 ? pht_3_128 : _GEN_3199; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3201 = 3'h3 == pht_windex & 8'h81 == _GEN_14976 ? pht_3_129 : _GEN_3200; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3202 = 3'h3 == pht_windex & 8'h82 == _GEN_14976 ? pht_3_130 : _GEN_3201; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3203 = 3'h3 == pht_windex & 8'h83 == _GEN_14976 ? pht_3_131 : _GEN_3202; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3204 = 3'h3 == pht_windex & 8'h84 == _GEN_14976 ? pht_3_132 : _GEN_3203; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3205 = 3'h3 == pht_windex & 8'h85 == _GEN_14976 ? pht_3_133 : _GEN_3204; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3206 = 3'h3 == pht_windex & 8'h86 == _GEN_14976 ? pht_3_134 : _GEN_3205; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3207 = 3'h3 == pht_windex & 8'h87 == _GEN_14976 ? pht_3_135 : _GEN_3206; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3208 = 3'h3 == pht_windex & 8'h88 == _GEN_14976 ? pht_3_136 : _GEN_3207; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3209 = 3'h3 == pht_windex & 8'h89 == _GEN_14976 ? pht_3_137 : _GEN_3208; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3210 = 3'h3 == pht_windex & 8'h8a == _GEN_14976 ? pht_3_138 : _GEN_3209; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3211 = 3'h3 == pht_windex & 8'h8b == _GEN_14976 ? pht_3_139 : _GEN_3210; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3212 = 3'h3 == pht_windex & 8'h8c == _GEN_14976 ? pht_3_140 : _GEN_3211; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3213 = 3'h3 == pht_windex & 8'h8d == _GEN_14976 ? pht_3_141 : _GEN_3212; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3214 = 3'h3 == pht_windex & 8'h8e == _GEN_14976 ? pht_3_142 : _GEN_3213; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3215 = 3'h3 == pht_windex & 8'h8f == _GEN_14976 ? pht_3_143 : _GEN_3214; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3216 = 3'h3 == pht_windex & 8'h90 == _GEN_14976 ? pht_3_144 : _GEN_3215; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3217 = 3'h3 == pht_windex & 8'h91 == _GEN_14976 ? pht_3_145 : _GEN_3216; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3218 = 3'h3 == pht_windex & 8'h92 == _GEN_14976 ? pht_3_146 : _GEN_3217; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3219 = 3'h3 == pht_windex & 8'h93 == _GEN_14976 ? pht_3_147 : _GEN_3218; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3220 = 3'h3 == pht_windex & 8'h94 == _GEN_14976 ? pht_3_148 : _GEN_3219; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3221 = 3'h3 == pht_windex & 8'h95 == _GEN_14976 ? pht_3_149 : _GEN_3220; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3222 = 3'h3 == pht_windex & 8'h96 == _GEN_14976 ? pht_3_150 : _GEN_3221; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3223 = 3'h3 == pht_windex & 8'h97 == _GEN_14976 ? pht_3_151 : _GEN_3222; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3224 = 3'h3 == pht_windex & 8'h98 == _GEN_14976 ? pht_3_152 : _GEN_3223; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3225 = 3'h3 == pht_windex & 8'h99 == _GEN_14976 ? pht_3_153 : _GEN_3224; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3226 = 3'h3 == pht_windex & 8'h9a == _GEN_14976 ? pht_3_154 : _GEN_3225; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3227 = 3'h3 == pht_windex & 8'h9b == _GEN_14976 ? pht_3_155 : _GEN_3226; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3228 = 3'h3 == pht_windex & 8'h9c == _GEN_14976 ? pht_3_156 : _GEN_3227; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3229 = 3'h3 == pht_windex & 8'h9d == _GEN_14976 ? pht_3_157 : _GEN_3228; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3230 = 3'h3 == pht_windex & 8'h9e == _GEN_14976 ? pht_3_158 : _GEN_3229; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3231 = 3'h3 == pht_windex & 8'h9f == _GEN_14976 ? pht_3_159 : _GEN_3230; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3232 = 3'h3 == pht_windex & 8'ha0 == _GEN_14976 ? pht_3_160 : _GEN_3231; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3233 = 3'h3 == pht_windex & 8'ha1 == _GEN_14976 ? pht_3_161 : _GEN_3232; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3234 = 3'h3 == pht_windex & 8'ha2 == _GEN_14976 ? pht_3_162 : _GEN_3233; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3235 = 3'h3 == pht_windex & 8'ha3 == _GEN_14976 ? pht_3_163 : _GEN_3234; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3236 = 3'h3 == pht_windex & 8'ha4 == _GEN_14976 ? pht_3_164 : _GEN_3235; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3237 = 3'h3 == pht_windex & 8'ha5 == _GEN_14976 ? pht_3_165 : _GEN_3236; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3238 = 3'h3 == pht_windex & 8'ha6 == _GEN_14976 ? pht_3_166 : _GEN_3237; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3239 = 3'h3 == pht_windex & 8'ha7 == _GEN_14976 ? pht_3_167 : _GEN_3238; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3240 = 3'h3 == pht_windex & 8'ha8 == _GEN_14976 ? pht_3_168 : _GEN_3239; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3241 = 3'h3 == pht_windex & 8'ha9 == _GEN_14976 ? pht_3_169 : _GEN_3240; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3242 = 3'h3 == pht_windex & 8'haa == _GEN_14976 ? pht_3_170 : _GEN_3241; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3243 = 3'h3 == pht_windex & 8'hab == _GEN_14976 ? pht_3_171 : _GEN_3242; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3244 = 3'h3 == pht_windex & 8'hac == _GEN_14976 ? pht_3_172 : _GEN_3243; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3245 = 3'h3 == pht_windex & 8'had == _GEN_14976 ? pht_3_173 : _GEN_3244; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3246 = 3'h3 == pht_windex & 8'hae == _GEN_14976 ? pht_3_174 : _GEN_3245; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3247 = 3'h3 == pht_windex & 8'haf == _GEN_14976 ? pht_3_175 : _GEN_3246; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3248 = 3'h3 == pht_windex & 8'hb0 == _GEN_14976 ? pht_3_176 : _GEN_3247; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3249 = 3'h3 == pht_windex & 8'hb1 == _GEN_14976 ? pht_3_177 : _GEN_3248; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3250 = 3'h3 == pht_windex & 8'hb2 == _GEN_14976 ? pht_3_178 : _GEN_3249; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3251 = 3'h3 == pht_windex & 8'hb3 == _GEN_14976 ? pht_3_179 : _GEN_3250; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3252 = 3'h3 == pht_windex & 8'hb4 == _GEN_14976 ? pht_3_180 : _GEN_3251; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3253 = 3'h3 == pht_windex & 8'hb5 == _GEN_14976 ? pht_3_181 : _GEN_3252; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3254 = 3'h3 == pht_windex & 8'hb6 == _GEN_14976 ? pht_3_182 : _GEN_3253; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3255 = 3'h3 == pht_windex & 8'hb7 == _GEN_14976 ? pht_3_183 : _GEN_3254; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3256 = 3'h3 == pht_windex & 8'hb8 == _GEN_14976 ? pht_3_184 : _GEN_3255; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3257 = 3'h3 == pht_windex & 8'hb9 == _GEN_14976 ? pht_3_185 : _GEN_3256; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3258 = 3'h3 == pht_windex & 8'hba == _GEN_14976 ? pht_3_186 : _GEN_3257; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3259 = 3'h3 == pht_windex & 8'hbb == _GEN_14976 ? pht_3_187 : _GEN_3258; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3260 = 3'h3 == pht_windex & 8'hbc == _GEN_14976 ? pht_3_188 : _GEN_3259; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3261 = 3'h3 == pht_windex & 8'hbd == _GEN_14976 ? pht_3_189 : _GEN_3260; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3262 = 3'h3 == pht_windex & 8'hbe == _GEN_14976 ? pht_3_190 : _GEN_3261; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3263 = 3'h3 == pht_windex & 8'hbf == _GEN_14976 ? pht_3_191 : _GEN_3262; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3264 = 3'h3 == pht_windex & 8'hc0 == _GEN_14976 ? pht_3_192 : _GEN_3263; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3265 = 3'h3 == pht_windex & 8'hc1 == _GEN_14976 ? pht_3_193 : _GEN_3264; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3266 = 3'h3 == pht_windex & 8'hc2 == _GEN_14976 ? pht_3_194 : _GEN_3265; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3267 = 3'h3 == pht_windex & 8'hc3 == _GEN_14976 ? pht_3_195 : _GEN_3266; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3268 = 3'h3 == pht_windex & 8'hc4 == _GEN_14976 ? pht_3_196 : _GEN_3267; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3269 = 3'h3 == pht_windex & 8'hc5 == _GEN_14976 ? pht_3_197 : _GEN_3268; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3270 = 3'h3 == pht_windex & 8'hc6 == _GEN_14976 ? pht_3_198 : _GEN_3269; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3271 = 3'h3 == pht_windex & 8'hc7 == _GEN_14976 ? pht_3_199 : _GEN_3270; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3272 = 3'h3 == pht_windex & 8'hc8 == _GEN_14976 ? pht_3_200 : _GEN_3271; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3273 = 3'h3 == pht_windex & 8'hc9 == _GEN_14976 ? pht_3_201 : _GEN_3272; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3274 = 3'h3 == pht_windex & 8'hca == _GEN_14976 ? pht_3_202 : _GEN_3273; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3275 = 3'h3 == pht_windex & 8'hcb == _GEN_14976 ? pht_3_203 : _GEN_3274; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3276 = 3'h3 == pht_windex & 8'hcc == _GEN_14976 ? pht_3_204 : _GEN_3275; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3277 = 3'h3 == pht_windex & 8'hcd == _GEN_14976 ? pht_3_205 : _GEN_3276; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3278 = 3'h3 == pht_windex & 8'hce == _GEN_14976 ? pht_3_206 : _GEN_3277; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3279 = 3'h3 == pht_windex & 8'hcf == _GEN_14976 ? pht_3_207 : _GEN_3278; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3280 = 3'h3 == pht_windex & 8'hd0 == _GEN_14976 ? pht_3_208 : _GEN_3279; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3281 = 3'h3 == pht_windex & 8'hd1 == _GEN_14976 ? pht_3_209 : _GEN_3280; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3282 = 3'h3 == pht_windex & 8'hd2 == _GEN_14976 ? pht_3_210 : _GEN_3281; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3283 = 3'h3 == pht_windex & 8'hd3 == _GEN_14976 ? pht_3_211 : _GEN_3282; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3284 = 3'h3 == pht_windex & 8'hd4 == _GEN_14976 ? pht_3_212 : _GEN_3283; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3285 = 3'h3 == pht_windex & 8'hd5 == _GEN_14976 ? pht_3_213 : _GEN_3284; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3286 = 3'h3 == pht_windex & 8'hd6 == _GEN_14976 ? pht_3_214 : _GEN_3285; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3287 = 3'h3 == pht_windex & 8'hd7 == _GEN_14976 ? pht_3_215 : _GEN_3286; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3288 = 3'h3 == pht_windex & 8'hd8 == _GEN_14976 ? pht_3_216 : _GEN_3287; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3289 = 3'h3 == pht_windex & 8'hd9 == _GEN_14976 ? pht_3_217 : _GEN_3288; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3290 = 3'h3 == pht_windex & 8'hda == _GEN_14976 ? pht_3_218 : _GEN_3289; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3291 = 3'h3 == pht_windex & 8'hdb == _GEN_14976 ? pht_3_219 : _GEN_3290; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3292 = 3'h3 == pht_windex & 8'hdc == _GEN_14976 ? pht_3_220 : _GEN_3291; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3293 = 3'h3 == pht_windex & 8'hdd == _GEN_14976 ? pht_3_221 : _GEN_3292; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3294 = 3'h3 == pht_windex & 8'hde == _GEN_14976 ? pht_3_222 : _GEN_3293; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3295 = 3'h3 == pht_windex & 8'hdf == _GEN_14976 ? pht_3_223 : _GEN_3294; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3296 = 3'h3 == pht_windex & 8'he0 == _GEN_14976 ? pht_3_224 : _GEN_3295; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3297 = 3'h3 == pht_windex & 8'he1 == _GEN_14976 ? pht_3_225 : _GEN_3296; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3298 = 3'h3 == pht_windex & 8'he2 == _GEN_14976 ? pht_3_226 : _GEN_3297; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3299 = 3'h3 == pht_windex & 8'he3 == _GEN_14976 ? pht_3_227 : _GEN_3298; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3300 = 3'h3 == pht_windex & 8'he4 == _GEN_14976 ? pht_3_228 : _GEN_3299; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3301 = 3'h3 == pht_windex & 8'he5 == _GEN_14976 ? pht_3_229 : _GEN_3300; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3302 = 3'h3 == pht_windex & 8'he6 == _GEN_14976 ? pht_3_230 : _GEN_3301; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3303 = 3'h3 == pht_windex & 8'he7 == _GEN_14976 ? pht_3_231 : _GEN_3302; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3304 = 3'h3 == pht_windex & 8'he8 == _GEN_14976 ? pht_3_232 : _GEN_3303; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3305 = 3'h3 == pht_windex & 8'he9 == _GEN_14976 ? pht_3_233 : _GEN_3304; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3306 = 3'h3 == pht_windex & 8'hea == _GEN_14976 ? pht_3_234 : _GEN_3305; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3307 = 3'h3 == pht_windex & 8'heb == _GEN_14976 ? pht_3_235 : _GEN_3306; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3308 = 3'h3 == pht_windex & 8'hec == _GEN_14976 ? pht_3_236 : _GEN_3307; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3309 = 3'h3 == pht_windex & 8'hed == _GEN_14976 ? pht_3_237 : _GEN_3308; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3310 = 3'h3 == pht_windex & 8'hee == _GEN_14976 ? pht_3_238 : _GEN_3309; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3311 = 3'h3 == pht_windex & 8'hef == _GEN_14976 ? pht_3_239 : _GEN_3310; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3312 = 3'h3 == pht_windex & 8'hf0 == _GEN_14976 ? pht_3_240 : _GEN_3311; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3313 = 3'h3 == pht_windex & 8'hf1 == _GEN_14976 ? pht_3_241 : _GEN_3312; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3314 = 3'h3 == pht_windex & 8'hf2 == _GEN_14976 ? pht_3_242 : _GEN_3313; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3315 = 3'h3 == pht_windex & 8'hf3 == _GEN_14976 ? pht_3_243 : _GEN_3314; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3316 = 3'h3 == pht_windex & 8'hf4 == _GEN_14976 ? pht_3_244 : _GEN_3315; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3317 = 3'h3 == pht_windex & 8'hf5 == _GEN_14976 ? pht_3_245 : _GEN_3316; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3318 = 3'h3 == pht_windex & 8'hf6 == _GEN_14976 ? pht_3_246 : _GEN_3317; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3319 = 3'h3 == pht_windex & 8'hf7 == _GEN_14976 ? pht_3_247 : _GEN_3318; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3320 = 3'h3 == pht_windex & 8'hf8 == _GEN_14976 ? pht_3_248 : _GEN_3319; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3321 = 3'h3 == pht_windex & 8'hf9 == _GEN_14976 ? pht_3_249 : _GEN_3320; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3322 = 3'h3 == pht_windex & 8'hfa == _GEN_14976 ? pht_3_250 : _GEN_3321; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3323 = 3'h3 == pht_windex & 8'hfb == _GEN_14976 ? pht_3_251 : _GEN_3322; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3324 = 3'h3 == pht_windex & 8'hfc == _GEN_14976 ? pht_3_252 : _GEN_3323; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3325 = 3'h3 == pht_windex & 8'hfd == _GEN_14976 ? pht_3_253 : _GEN_3324; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3326 = 3'h3 == pht_windex & 8'hfe == _GEN_14976 ? pht_3_254 : _GEN_3325; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3327 = 3'h3 == pht_windex & 8'hff == _GEN_14976 ? pht_3_255 : _GEN_3326; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_17472 = 3'h4 == pht_windex; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3328 = 3'h4 == pht_windex & 6'h0 == pht_waddr ? pht_4_0 : _GEN_3327; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3329 = 3'h4 == pht_windex & 6'h1 == pht_waddr ? pht_4_1 : _GEN_3328; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3330 = 3'h4 == pht_windex & 6'h2 == pht_waddr ? pht_4_2 : _GEN_3329; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3331 = 3'h4 == pht_windex & 6'h3 == pht_waddr ? pht_4_3 : _GEN_3330; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3332 = 3'h4 == pht_windex & 6'h4 == pht_waddr ? pht_4_4 : _GEN_3331; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3333 = 3'h4 == pht_windex & 6'h5 == pht_waddr ? pht_4_5 : _GEN_3332; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3334 = 3'h4 == pht_windex & 6'h6 == pht_waddr ? pht_4_6 : _GEN_3333; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3335 = 3'h4 == pht_windex & 6'h7 == pht_waddr ? pht_4_7 : _GEN_3334; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3336 = 3'h4 == pht_windex & 6'h8 == pht_waddr ? pht_4_8 : _GEN_3335; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3337 = 3'h4 == pht_windex & 6'h9 == pht_waddr ? pht_4_9 : _GEN_3336; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3338 = 3'h4 == pht_windex & 6'ha == pht_waddr ? pht_4_10 : _GEN_3337; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3339 = 3'h4 == pht_windex & 6'hb == pht_waddr ? pht_4_11 : _GEN_3338; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3340 = 3'h4 == pht_windex & 6'hc == pht_waddr ? pht_4_12 : _GEN_3339; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3341 = 3'h4 == pht_windex & 6'hd == pht_waddr ? pht_4_13 : _GEN_3340; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3342 = 3'h4 == pht_windex & 6'he == pht_waddr ? pht_4_14 : _GEN_3341; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3343 = 3'h4 == pht_windex & 6'hf == pht_waddr ? pht_4_15 : _GEN_3342; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3344 = 3'h4 == pht_windex & 6'h10 == pht_waddr ? pht_4_16 : _GEN_3343; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3345 = 3'h4 == pht_windex & 6'h11 == pht_waddr ? pht_4_17 : _GEN_3344; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3346 = 3'h4 == pht_windex & 6'h12 == pht_waddr ? pht_4_18 : _GEN_3345; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3347 = 3'h4 == pht_windex & 6'h13 == pht_waddr ? pht_4_19 : _GEN_3346; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3348 = 3'h4 == pht_windex & 6'h14 == pht_waddr ? pht_4_20 : _GEN_3347; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3349 = 3'h4 == pht_windex & 6'h15 == pht_waddr ? pht_4_21 : _GEN_3348; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3350 = 3'h4 == pht_windex & 6'h16 == pht_waddr ? pht_4_22 : _GEN_3349; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3351 = 3'h4 == pht_windex & 6'h17 == pht_waddr ? pht_4_23 : _GEN_3350; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3352 = 3'h4 == pht_windex & 6'h18 == pht_waddr ? pht_4_24 : _GEN_3351; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3353 = 3'h4 == pht_windex & 6'h19 == pht_waddr ? pht_4_25 : _GEN_3352; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3354 = 3'h4 == pht_windex & 6'h1a == pht_waddr ? pht_4_26 : _GEN_3353; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3355 = 3'h4 == pht_windex & 6'h1b == pht_waddr ? pht_4_27 : _GEN_3354; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3356 = 3'h4 == pht_windex & 6'h1c == pht_waddr ? pht_4_28 : _GEN_3355; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3357 = 3'h4 == pht_windex & 6'h1d == pht_waddr ? pht_4_29 : _GEN_3356; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3358 = 3'h4 == pht_windex & 6'h1e == pht_waddr ? pht_4_30 : _GEN_3357; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3359 = 3'h4 == pht_windex & 6'h1f == pht_waddr ? pht_4_31 : _GEN_3358; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3360 = 3'h4 == pht_windex & 6'h20 == pht_waddr ? pht_4_32 : _GEN_3359; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3361 = 3'h4 == pht_windex & 6'h21 == pht_waddr ? pht_4_33 : _GEN_3360; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3362 = 3'h4 == pht_windex & 6'h22 == pht_waddr ? pht_4_34 : _GEN_3361; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3363 = 3'h4 == pht_windex & 6'h23 == pht_waddr ? pht_4_35 : _GEN_3362; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3364 = 3'h4 == pht_windex & 6'h24 == pht_waddr ? pht_4_36 : _GEN_3363; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3365 = 3'h4 == pht_windex & 6'h25 == pht_waddr ? pht_4_37 : _GEN_3364; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3366 = 3'h4 == pht_windex & 6'h26 == pht_waddr ? pht_4_38 : _GEN_3365; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3367 = 3'h4 == pht_windex & 6'h27 == pht_waddr ? pht_4_39 : _GEN_3366; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3368 = 3'h4 == pht_windex & 6'h28 == pht_waddr ? pht_4_40 : _GEN_3367; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3369 = 3'h4 == pht_windex & 6'h29 == pht_waddr ? pht_4_41 : _GEN_3368; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3370 = 3'h4 == pht_windex & 6'h2a == pht_waddr ? pht_4_42 : _GEN_3369; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3371 = 3'h4 == pht_windex & 6'h2b == pht_waddr ? pht_4_43 : _GEN_3370; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3372 = 3'h4 == pht_windex & 6'h2c == pht_waddr ? pht_4_44 : _GEN_3371; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3373 = 3'h4 == pht_windex & 6'h2d == pht_waddr ? pht_4_45 : _GEN_3372; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3374 = 3'h4 == pht_windex & 6'h2e == pht_waddr ? pht_4_46 : _GEN_3373; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3375 = 3'h4 == pht_windex & 6'h2f == pht_waddr ? pht_4_47 : _GEN_3374; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3376 = 3'h4 == pht_windex & 6'h30 == pht_waddr ? pht_4_48 : _GEN_3375; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3377 = 3'h4 == pht_windex & 6'h31 == pht_waddr ? pht_4_49 : _GEN_3376; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3378 = 3'h4 == pht_windex & 6'h32 == pht_waddr ? pht_4_50 : _GEN_3377; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3379 = 3'h4 == pht_windex & 6'h33 == pht_waddr ? pht_4_51 : _GEN_3378; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3380 = 3'h4 == pht_windex & 6'h34 == pht_waddr ? pht_4_52 : _GEN_3379; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3381 = 3'h4 == pht_windex & 6'h35 == pht_waddr ? pht_4_53 : _GEN_3380; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3382 = 3'h4 == pht_windex & 6'h36 == pht_waddr ? pht_4_54 : _GEN_3381; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3383 = 3'h4 == pht_windex & 6'h37 == pht_waddr ? pht_4_55 : _GEN_3382; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3384 = 3'h4 == pht_windex & 6'h38 == pht_waddr ? pht_4_56 : _GEN_3383; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3385 = 3'h4 == pht_windex & 6'h39 == pht_waddr ? pht_4_57 : _GEN_3384; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3386 = 3'h4 == pht_windex & 6'h3a == pht_waddr ? pht_4_58 : _GEN_3385; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3387 = 3'h4 == pht_windex & 6'h3b == pht_waddr ? pht_4_59 : _GEN_3386; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3388 = 3'h4 == pht_windex & 6'h3c == pht_waddr ? pht_4_60 : _GEN_3387; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3389 = 3'h4 == pht_windex & 6'h3d == pht_waddr ? pht_4_61 : _GEN_3388; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3390 = 3'h4 == pht_windex & 6'h3e == pht_waddr ? pht_4_62 : _GEN_3389; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3391 = 3'h4 == pht_windex & 6'h3f == pht_waddr ? pht_4_63 : _GEN_3390; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3392 = 3'h4 == pht_windex & 7'h40 == _GEN_14784 ? pht_4_64 : _GEN_3391; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3393 = 3'h4 == pht_windex & 7'h41 == _GEN_14784 ? pht_4_65 : _GEN_3392; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3394 = 3'h4 == pht_windex & 7'h42 == _GEN_14784 ? pht_4_66 : _GEN_3393; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3395 = 3'h4 == pht_windex & 7'h43 == _GEN_14784 ? pht_4_67 : _GEN_3394; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3396 = 3'h4 == pht_windex & 7'h44 == _GEN_14784 ? pht_4_68 : _GEN_3395; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3397 = 3'h4 == pht_windex & 7'h45 == _GEN_14784 ? pht_4_69 : _GEN_3396; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3398 = 3'h4 == pht_windex & 7'h46 == _GEN_14784 ? pht_4_70 : _GEN_3397; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3399 = 3'h4 == pht_windex & 7'h47 == _GEN_14784 ? pht_4_71 : _GEN_3398; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3400 = 3'h4 == pht_windex & 7'h48 == _GEN_14784 ? pht_4_72 : _GEN_3399; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3401 = 3'h4 == pht_windex & 7'h49 == _GEN_14784 ? pht_4_73 : _GEN_3400; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3402 = 3'h4 == pht_windex & 7'h4a == _GEN_14784 ? pht_4_74 : _GEN_3401; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3403 = 3'h4 == pht_windex & 7'h4b == _GEN_14784 ? pht_4_75 : _GEN_3402; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3404 = 3'h4 == pht_windex & 7'h4c == _GEN_14784 ? pht_4_76 : _GEN_3403; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3405 = 3'h4 == pht_windex & 7'h4d == _GEN_14784 ? pht_4_77 : _GEN_3404; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3406 = 3'h4 == pht_windex & 7'h4e == _GEN_14784 ? pht_4_78 : _GEN_3405; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3407 = 3'h4 == pht_windex & 7'h4f == _GEN_14784 ? pht_4_79 : _GEN_3406; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3408 = 3'h4 == pht_windex & 7'h50 == _GEN_14784 ? pht_4_80 : _GEN_3407; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3409 = 3'h4 == pht_windex & 7'h51 == _GEN_14784 ? pht_4_81 : _GEN_3408; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3410 = 3'h4 == pht_windex & 7'h52 == _GEN_14784 ? pht_4_82 : _GEN_3409; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3411 = 3'h4 == pht_windex & 7'h53 == _GEN_14784 ? pht_4_83 : _GEN_3410; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3412 = 3'h4 == pht_windex & 7'h54 == _GEN_14784 ? pht_4_84 : _GEN_3411; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3413 = 3'h4 == pht_windex & 7'h55 == _GEN_14784 ? pht_4_85 : _GEN_3412; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3414 = 3'h4 == pht_windex & 7'h56 == _GEN_14784 ? pht_4_86 : _GEN_3413; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3415 = 3'h4 == pht_windex & 7'h57 == _GEN_14784 ? pht_4_87 : _GEN_3414; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3416 = 3'h4 == pht_windex & 7'h58 == _GEN_14784 ? pht_4_88 : _GEN_3415; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3417 = 3'h4 == pht_windex & 7'h59 == _GEN_14784 ? pht_4_89 : _GEN_3416; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3418 = 3'h4 == pht_windex & 7'h5a == _GEN_14784 ? pht_4_90 : _GEN_3417; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3419 = 3'h4 == pht_windex & 7'h5b == _GEN_14784 ? pht_4_91 : _GEN_3418; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3420 = 3'h4 == pht_windex & 7'h5c == _GEN_14784 ? pht_4_92 : _GEN_3419; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3421 = 3'h4 == pht_windex & 7'h5d == _GEN_14784 ? pht_4_93 : _GEN_3420; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3422 = 3'h4 == pht_windex & 7'h5e == _GEN_14784 ? pht_4_94 : _GEN_3421; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3423 = 3'h4 == pht_windex & 7'h5f == _GEN_14784 ? pht_4_95 : _GEN_3422; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3424 = 3'h4 == pht_windex & 7'h60 == _GEN_14784 ? pht_4_96 : _GEN_3423; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3425 = 3'h4 == pht_windex & 7'h61 == _GEN_14784 ? pht_4_97 : _GEN_3424; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3426 = 3'h4 == pht_windex & 7'h62 == _GEN_14784 ? pht_4_98 : _GEN_3425; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3427 = 3'h4 == pht_windex & 7'h63 == _GEN_14784 ? pht_4_99 : _GEN_3426; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3428 = 3'h4 == pht_windex & 7'h64 == _GEN_14784 ? pht_4_100 : _GEN_3427; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3429 = 3'h4 == pht_windex & 7'h65 == _GEN_14784 ? pht_4_101 : _GEN_3428; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3430 = 3'h4 == pht_windex & 7'h66 == _GEN_14784 ? pht_4_102 : _GEN_3429; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3431 = 3'h4 == pht_windex & 7'h67 == _GEN_14784 ? pht_4_103 : _GEN_3430; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3432 = 3'h4 == pht_windex & 7'h68 == _GEN_14784 ? pht_4_104 : _GEN_3431; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3433 = 3'h4 == pht_windex & 7'h69 == _GEN_14784 ? pht_4_105 : _GEN_3432; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3434 = 3'h4 == pht_windex & 7'h6a == _GEN_14784 ? pht_4_106 : _GEN_3433; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3435 = 3'h4 == pht_windex & 7'h6b == _GEN_14784 ? pht_4_107 : _GEN_3434; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3436 = 3'h4 == pht_windex & 7'h6c == _GEN_14784 ? pht_4_108 : _GEN_3435; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3437 = 3'h4 == pht_windex & 7'h6d == _GEN_14784 ? pht_4_109 : _GEN_3436; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3438 = 3'h4 == pht_windex & 7'h6e == _GEN_14784 ? pht_4_110 : _GEN_3437; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3439 = 3'h4 == pht_windex & 7'h6f == _GEN_14784 ? pht_4_111 : _GEN_3438; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3440 = 3'h4 == pht_windex & 7'h70 == _GEN_14784 ? pht_4_112 : _GEN_3439; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3441 = 3'h4 == pht_windex & 7'h71 == _GEN_14784 ? pht_4_113 : _GEN_3440; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3442 = 3'h4 == pht_windex & 7'h72 == _GEN_14784 ? pht_4_114 : _GEN_3441; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3443 = 3'h4 == pht_windex & 7'h73 == _GEN_14784 ? pht_4_115 : _GEN_3442; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3444 = 3'h4 == pht_windex & 7'h74 == _GEN_14784 ? pht_4_116 : _GEN_3443; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3445 = 3'h4 == pht_windex & 7'h75 == _GEN_14784 ? pht_4_117 : _GEN_3444; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3446 = 3'h4 == pht_windex & 7'h76 == _GEN_14784 ? pht_4_118 : _GEN_3445; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3447 = 3'h4 == pht_windex & 7'h77 == _GEN_14784 ? pht_4_119 : _GEN_3446; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3448 = 3'h4 == pht_windex & 7'h78 == _GEN_14784 ? pht_4_120 : _GEN_3447; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3449 = 3'h4 == pht_windex & 7'h79 == _GEN_14784 ? pht_4_121 : _GEN_3448; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3450 = 3'h4 == pht_windex & 7'h7a == _GEN_14784 ? pht_4_122 : _GEN_3449; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3451 = 3'h4 == pht_windex & 7'h7b == _GEN_14784 ? pht_4_123 : _GEN_3450; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3452 = 3'h4 == pht_windex & 7'h7c == _GEN_14784 ? pht_4_124 : _GEN_3451; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3453 = 3'h4 == pht_windex & 7'h7d == _GEN_14784 ? pht_4_125 : _GEN_3452; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3454 = 3'h4 == pht_windex & 7'h7e == _GEN_14784 ? pht_4_126 : _GEN_3453; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3455 = 3'h4 == pht_windex & 7'h7f == _GEN_14784 ? pht_4_127 : _GEN_3454; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3456 = 3'h4 == pht_windex & 8'h80 == _GEN_14976 ? pht_4_128 : _GEN_3455; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3457 = 3'h4 == pht_windex & 8'h81 == _GEN_14976 ? pht_4_129 : _GEN_3456; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3458 = 3'h4 == pht_windex & 8'h82 == _GEN_14976 ? pht_4_130 : _GEN_3457; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3459 = 3'h4 == pht_windex & 8'h83 == _GEN_14976 ? pht_4_131 : _GEN_3458; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3460 = 3'h4 == pht_windex & 8'h84 == _GEN_14976 ? pht_4_132 : _GEN_3459; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3461 = 3'h4 == pht_windex & 8'h85 == _GEN_14976 ? pht_4_133 : _GEN_3460; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3462 = 3'h4 == pht_windex & 8'h86 == _GEN_14976 ? pht_4_134 : _GEN_3461; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3463 = 3'h4 == pht_windex & 8'h87 == _GEN_14976 ? pht_4_135 : _GEN_3462; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3464 = 3'h4 == pht_windex & 8'h88 == _GEN_14976 ? pht_4_136 : _GEN_3463; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3465 = 3'h4 == pht_windex & 8'h89 == _GEN_14976 ? pht_4_137 : _GEN_3464; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3466 = 3'h4 == pht_windex & 8'h8a == _GEN_14976 ? pht_4_138 : _GEN_3465; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3467 = 3'h4 == pht_windex & 8'h8b == _GEN_14976 ? pht_4_139 : _GEN_3466; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3468 = 3'h4 == pht_windex & 8'h8c == _GEN_14976 ? pht_4_140 : _GEN_3467; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3469 = 3'h4 == pht_windex & 8'h8d == _GEN_14976 ? pht_4_141 : _GEN_3468; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3470 = 3'h4 == pht_windex & 8'h8e == _GEN_14976 ? pht_4_142 : _GEN_3469; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3471 = 3'h4 == pht_windex & 8'h8f == _GEN_14976 ? pht_4_143 : _GEN_3470; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3472 = 3'h4 == pht_windex & 8'h90 == _GEN_14976 ? pht_4_144 : _GEN_3471; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3473 = 3'h4 == pht_windex & 8'h91 == _GEN_14976 ? pht_4_145 : _GEN_3472; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3474 = 3'h4 == pht_windex & 8'h92 == _GEN_14976 ? pht_4_146 : _GEN_3473; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3475 = 3'h4 == pht_windex & 8'h93 == _GEN_14976 ? pht_4_147 : _GEN_3474; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3476 = 3'h4 == pht_windex & 8'h94 == _GEN_14976 ? pht_4_148 : _GEN_3475; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3477 = 3'h4 == pht_windex & 8'h95 == _GEN_14976 ? pht_4_149 : _GEN_3476; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3478 = 3'h4 == pht_windex & 8'h96 == _GEN_14976 ? pht_4_150 : _GEN_3477; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3479 = 3'h4 == pht_windex & 8'h97 == _GEN_14976 ? pht_4_151 : _GEN_3478; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3480 = 3'h4 == pht_windex & 8'h98 == _GEN_14976 ? pht_4_152 : _GEN_3479; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3481 = 3'h4 == pht_windex & 8'h99 == _GEN_14976 ? pht_4_153 : _GEN_3480; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3482 = 3'h4 == pht_windex & 8'h9a == _GEN_14976 ? pht_4_154 : _GEN_3481; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3483 = 3'h4 == pht_windex & 8'h9b == _GEN_14976 ? pht_4_155 : _GEN_3482; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3484 = 3'h4 == pht_windex & 8'h9c == _GEN_14976 ? pht_4_156 : _GEN_3483; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3485 = 3'h4 == pht_windex & 8'h9d == _GEN_14976 ? pht_4_157 : _GEN_3484; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3486 = 3'h4 == pht_windex & 8'h9e == _GEN_14976 ? pht_4_158 : _GEN_3485; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3487 = 3'h4 == pht_windex & 8'h9f == _GEN_14976 ? pht_4_159 : _GEN_3486; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3488 = 3'h4 == pht_windex & 8'ha0 == _GEN_14976 ? pht_4_160 : _GEN_3487; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3489 = 3'h4 == pht_windex & 8'ha1 == _GEN_14976 ? pht_4_161 : _GEN_3488; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3490 = 3'h4 == pht_windex & 8'ha2 == _GEN_14976 ? pht_4_162 : _GEN_3489; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3491 = 3'h4 == pht_windex & 8'ha3 == _GEN_14976 ? pht_4_163 : _GEN_3490; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3492 = 3'h4 == pht_windex & 8'ha4 == _GEN_14976 ? pht_4_164 : _GEN_3491; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3493 = 3'h4 == pht_windex & 8'ha5 == _GEN_14976 ? pht_4_165 : _GEN_3492; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3494 = 3'h4 == pht_windex & 8'ha6 == _GEN_14976 ? pht_4_166 : _GEN_3493; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3495 = 3'h4 == pht_windex & 8'ha7 == _GEN_14976 ? pht_4_167 : _GEN_3494; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3496 = 3'h4 == pht_windex & 8'ha8 == _GEN_14976 ? pht_4_168 : _GEN_3495; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3497 = 3'h4 == pht_windex & 8'ha9 == _GEN_14976 ? pht_4_169 : _GEN_3496; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3498 = 3'h4 == pht_windex & 8'haa == _GEN_14976 ? pht_4_170 : _GEN_3497; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3499 = 3'h4 == pht_windex & 8'hab == _GEN_14976 ? pht_4_171 : _GEN_3498; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3500 = 3'h4 == pht_windex & 8'hac == _GEN_14976 ? pht_4_172 : _GEN_3499; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3501 = 3'h4 == pht_windex & 8'had == _GEN_14976 ? pht_4_173 : _GEN_3500; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3502 = 3'h4 == pht_windex & 8'hae == _GEN_14976 ? pht_4_174 : _GEN_3501; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3503 = 3'h4 == pht_windex & 8'haf == _GEN_14976 ? pht_4_175 : _GEN_3502; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3504 = 3'h4 == pht_windex & 8'hb0 == _GEN_14976 ? pht_4_176 : _GEN_3503; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3505 = 3'h4 == pht_windex & 8'hb1 == _GEN_14976 ? pht_4_177 : _GEN_3504; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3506 = 3'h4 == pht_windex & 8'hb2 == _GEN_14976 ? pht_4_178 : _GEN_3505; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3507 = 3'h4 == pht_windex & 8'hb3 == _GEN_14976 ? pht_4_179 : _GEN_3506; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3508 = 3'h4 == pht_windex & 8'hb4 == _GEN_14976 ? pht_4_180 : _GEN_3507; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3509 = 3'h4 == pht_windex & 8'hb5 == _GEN_14976 ? pht_4_181 : _GEN_3508; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3510 = 3'h4 == pht_windex & 8'hb6 == _GEN_14976 ? pht_4_182 : _GEN_3509; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3511 = 3'h4 == pht_windex & 8'hb7 == _GEN_14976 ? pht_4_183 : _GEN_3510; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3512 = 3'h4 == pht_windex & 8'hb8 == _GEN_14976 ? pht_4_184 : _GEN_3511; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3513 = 3'h4 == pht_windex & 8'hb9 == _GEN_14976 ? pht_4_185 : _GEN_3512; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3514 = 3'h4 == pht_windex & 8'hba == _GEN_14976 ? pht_4_186 : _GEN_3513; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3515 = 3'h4 == pht_windex & 8'hbb == _GEN_14976 ? pht_4_187 : _GEN_3514; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3516 = 3'h4 == pht_windex & 8'hbc == _GEN_14976 ? pht_4_188 : _GEN_3515; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3517 = 3'h4 == pht_windex & 8'hbd == _GEN_14976 ? pht_4_189 : _GEN_3516; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3518 = 3'h4 == pht_windex & 8'hbe == _GEN_14976 ? pht_4_190 : _GEN_3517; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3519 = 3'h4 == pht_windex & 8'hbf == _GEN_14976 ? pht_4_191 : _GEN_3518; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3520 = 3'h4 == pht_windex & 8'hc0 == _GEN_14976 ? pht_4_192 : _GEN_3519; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3521 = 3'h4 == pht_windex & 8'hc1 == _GEN_14976 ? pht_4_193 : _GEN_3520; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3522 = 3'h4 == pht_windex & 8'hc2 == _GEN_14976 ? pht_4_194 : _GEN_3521; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3523 = 3'h4 == pht_windex & 8'hc3 == _GEN_14976 ? pht_4_195 : _GEN_3522; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3524 = 3'h4 == pht_windex & 8'hc4 == _GEN_14976 ? pht_4_196 : _GEN_3523; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3525 = 3'h4 == pht_windex & 8'hc5 == _GEN_14976 ? pht_4_197 : _GEN_3524; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3526 = 3'h4 == pht_windex & 8'hc6 == _GEN_14976 ? pht_4_198 : _GEN_3525; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3527 = 3'h4 == pht_windex & 8'hc7 == _GEN_14976 ? pht_4_199 : _GEN_3526; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3528 = 3'h4 == pht_windex & 8'hc8 == _GEN_14976 ? pht_4_200 : _GEN_3527; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3529 = 3'h4 == pht_windex & 8'hc9 == _GEN_14976 ? pht_4_201 : _GEN_3528; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3530 = 3'h4 == pht_windex & 8'hca == _GEN_14976 ? pht_4_202 : _GEN_3529; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3531 = 3'h4 == pht_windex & 8'hcb == _GEN_14976 ? pht_4_203 : _GEN_3530; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3532 = 3'h4 == pht_windex & 8'hcc == _GEN_14976 ? pht_4_204 : _GEN_3531; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3533 = 3'h4 == pht_windex & 8'hcd == _GEN_14976 ? pht_4_205 : _GEN_3532; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3534 = 3'h4 == pht_windex & 8'hce == _GEN_14976 ? pht_4_206 : _GEN_3533; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3535 = 3'h4 == pht_windex & 8'hcf == _GEN_14976 ? pht_4_207 : _GEN_3534; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3536 = 3'h4 == pht_windex & 8'hd0 == _GEN_14976 ? pht_4_208 : _GEN_3535; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3537 = 3'h4 == pht_windex & 8'hd1 == _GEN_14976 ? pht_4_209 : _GEN_3536; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3538 = 3'h4 == pht_windex & 8'hd2 == _GEN_14976 ? pht_4_210 : _GEN_3537; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3539 = 3'h4 == pht_windex & 8'hd3 == _GEN_14976 ? pht_4_211 : _GEN_3538; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3540 = 3'h4 == pht_windex & 8'hd4 == _GEN_14976 ? pht_4_212 : _GEN_3539; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3541 = 3'h4 == pht_windex & 8'hd5 == _GEN_14976 ? pht_4_213 : _GEN_3540; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3542 = 3'h4 == pht_windex & 8'hd6 == _GEN_14976 ? pht_4_214 : _GEN_3541; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3543 = 3'h4 == pht_windex & 8'hd7 == _GEN_14976 ? pht_4_215 : _GEN_3542; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3544 = 3'h4 == pht_windex & 8'hd8 == _GEN_14976 ? pht_4_216 : _GEN_3543; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3545 = 3'h4 == pht_windex & 8'hd9 == _GEN_14976 ? pht_4_217 : _GEN_3544; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3546 = 3'h4 == pht_windex & 8'hda == _GEN_14976 ? pht_4_218 : _GEN_3545; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3547 = 3'h4 == pht_windex & 8'hdb == _GEN_14976 ? pht_4_219 : _GEN_3546; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3548 = 3'h4 == pht_windex & 8'hdc == _GEN_14976 ? pht_4_220 : _GEN_3547; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3549 = 3'h4 == pht_windex & 8'hdd == _GEN_14976 ? pht_4_221 : _GEN_3548; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3550 = 3'h4 == pht_windex & 8'hde == _GEN_14976 ? pht_4_222 : _GEN_3549; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3551 = 3'h4 == pht_windex & 8'hdf == _GEN_14976 ? pht_4_223 : _GEN_3550; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3552 = 3'h4 == pht_windex & 8'he0 == _GEN_14976 ? pht_4_224 : _GEN_3551; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3553 = 3'h4 == pht_windex & 8'he1 == _GEN_14976 ? pht_4_225 : _GEN_3552; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3554 = 3'h4 == pht_windex & 8'he2 == _GEN_14976 ? pht_4_226 : _GEN_3553; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3555 = 3'h4 == pht_windex & 8'he3 == _GEN_14976 ? pht_4_227 : _GEN_3554; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3556 = 3'h4 == pht_windex & 8'he4 == _GEN_14976 ? pht_4_228 : _GEN_3555; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3557 = 3'h4 == pht_windex & 8'he5 == _GEN_14976 ? pht_4_229 : _GEN_3556; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3558 = 3'h4 == pht_windex & 8'he6 == _GEN_14976 ? pht_4_230 : _GEN_3557; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3559 = 3'h4 == pht_windex & 8'he7 == _GEN_14976 ? pht_4_231 : _GEN_3558; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3560 = 3'h4 == pht_windex & 8'he8 == _GEN_14976 ? pht_4_232 : _GEN_3559; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3561 = 3'h4 == pht_windex & 8'he9 == _GEN_14976 ? pht_4_233 : _GEN_3560; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3562 = 3'h4 == pht_windex & 8'hea == _GEN_14976 ? pht_4_234 : _GEN_3561; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3563 = 3'h4 == pht_windex & 8'heb == _GEN_14976 ? pht_4_235 : _GEN_3562; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3564 = 3'h4 == pht_windex & 8'hec == _GEN_14976 ? pht_4_236 : _GEN_3563; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3565 = 3'h4 == pht_windex & 8'hed == _GEN_14976 ? pht_4_237 : _GEN_3564; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3566 = 3'h4 == pht_windex & 8'hee == _GEN_14976 ? pht_4_238 : _GEN_3565; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3567 = 3'h4 == pht_windex & 8'hef == _GEN_14976 ? pht_4_239 : _GEN_3566; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3568 = 3'h4 == pht_windex & 8'hf0 == _GEN_14976 ? pht_4_240 : _GEN_3567; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3569 = 3'h4 == pht_windex & 8'hf1 == _GEN_14976 ? pht_4_241 : _GEN_3568; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3570 = 3'h4 == pht_windex & 8'hf2 == _GEN_14976 ? pht_4_242 : _GEN_3569; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3571 = 3'h4 == pht_windex & 8'hf3 == _GEN_14976 ? pht_4_243 : _GEN_3570; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3572 = 3'h4 == pht_windex & 8'hf4 == _GEN_14976 ? pht_4_244 : _GEN_3571; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3573 = 3'h4 == pht_windex & 8'hf5 == _GEN_14976 ? pht_4_245 : _GEN_3572; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3574 = 3'h4 == pht_windex & 8'hf6 == _GEN_14976 ? pht_4_246 : _GEN_3573; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3575 = 3'h4 == pht_windex & 8'hf7 == _GEN_14976 ? pht_4_247 : _GEN_3574; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3576 = 3'h4 == pht_windex & 8'hf8 == _GEN_14976 ? pht_4_248 : _GEN_3575; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3577 = 3'h4 == pht_windex & 8'hf9 == _GEN_14976 ? pht_4_249 : _GEN_3576; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3578 = 3'h4 == pht_windex & 8'hfa == _GEN_14976 ? pht_4_250 : _GEN_3577; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3579 = 3'h4 == pht_windex & 8'hfb == _GEN_14976 ? pht_4_251 : _GEN_3578; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3580 = 3'h4 == pht_windex & 8'hfc == _GEN_14976 ? pht_4_252 : _GEN_3579; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3581 = 3'h4 == pht_windex & 8'hfd == _GEN_14976 ? pht_4_253 : _GEN_3580; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3582 = 3'h4 == pht_windex & 8'hfe == _GEN_14976 ? pht_4_254 : _GEN_3581; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3583 = 3'h4 == pht_windex & 8'hff == _GEN_14976 ? pht_4_255 : _GEN_3582; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_18176 = 3'h5 == pht_windex; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3584 = 3'h5 == pht_windex & 6'h0 == pht_waddr ? pht_5_0 : _GEN_3583; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3585 = 3'h5 == pht_windex & 6'h1 == pht_waddr ? pht_5_1 : _GEN_3584; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3586 = 3'h5 == pht_windex & 6'h2 == pht_waddr ? pht_5_2 : _GEN_3585; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3587 = 3'h5 == pht_windex & 6'h3 == pht_waddr ? pht_5_3 : _GEN_3586; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3588 = 3'h5 == pht_windex & 6'h4 == pht_waddr ? pht_5_4 : _GEN_3587; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3589 = 3'h5 == pht_windex & 6'h5 == pht_waddr ? pht_5_5 : _GEN_3588; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3590 = 3'h5 == pht_windex & 6'h6 == pht_waddr ? pht_5_6 : _GEN_3589; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3591 = 3'h5 == pht_windex & 6'h7 == pht_waddr ? pht_5_7 : _GEN_3590; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3592 = 3'h5 == pht_windex & 6'h8 == pht_waddr ? pht_5_8 : _GEN_3591; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3593 = 3'h5 == pht_windex & 6'h9 == pht_waddr ? pht_5_9 : _GEN_3592; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3594 = 3'h5 == pht_windex & 6'ha == pht_waddr ? pht_5_10 : _GEN_3593; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3595 = 3'h5 == pht_windex & 6'hb == pht_waddr ? pht_5_11 : _GEN_3594; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3596 = 3'h5 == pht_windex & 6'hc == pht_waddr ? pht_5_12 : _GEN_3595; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3597 = 3'h5 == pht_windex & 6'hd == pht_waddr ? pht_5_13 : _GEN_3596; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3598 = 3'h5 == pht_windex & 6'he == pht_waddr ? pht_5_14 : _GEN_3597; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3599 = 3'h5 == pht_windex & 6'hf == pht_waddr ? pht_5_15 : _GEN_3598; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3600 = 3'h5 == pht_windex & 6'h10 == pht_waddr ? pht_5_16 : _GEN_3599; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3601 = 3'h5 == pht_windex & 6'h11 == pht_waddr ? pht_5_17 : _GEN_3600; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3602 = 3'h5 == pht_windex & 6'h12 == pht_waddr ? pht_5_18 : _GEN_3601; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3603 = 3'h5 == pht_windex & 6'h13 == pht_waddr ? pht_5_19 : _GEN_3602; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3604 = 3'h5 == pht_windex & 6'h14 == pht_waddr ? pht_5_20 : _GEN_3603; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3605 = 3'h5 == pht_windex & 6'h15 == pht_waddr ? pht_5_21 : _GEN_3604; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3606 = 3'h5 == pht_windex & 6'h16 == pht_waddr ? pht_5_22 : _GEN_3605; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3607 = 3'h5 == pht_windex & 6'h17 == pht_waddr ? pht_5_23 : _GEN_3606; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3608 = 3'h5 == pht_windex & 6'h18 == pht_waddr ? pht_5_24 : _GEN_3607; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3609 = 3'h5 == pht_windex & 6'h19 == pht_waddr ? pht_5_25 : _GEN_3608; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3610 = 3'h5 == pht_windex & 6'h1a == pht_waddr ? pht_5_26 : _GEN_3609; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3611 = 3'h5 == pht_windex & 6'h1b == pht_waddr ? pht_5_27 : _GEN_3610; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3612 = 3'h5 == pht_windex & 6'h1c == pht_waddr ? pht_5_28 : _GEN_3611; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3613 = 3'h5 == pht_windex & 6'h1d == pht_waddr ? pht_5_29 : _GEN_3612; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3614 = 3'h5 == pht_windex & 6'h1e == pht_waddr ? pht_5_30 : _GEN_3613; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3615 = 3'h5 == pht_windex & 6'h1f == pht_waddr ? pht_5_31 : _GEN_3614; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3616 = 3'h5 == pht_windex & 6'h20 == pht_waddr ? pht_5_32 : _GEN_3615; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3617 = 3'h5 == pht_windex & 6'h21 == pht_waddr ? pht_5_33 : _GEN_3616; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3618 = 3'h5 == pht_windex & 6'h22 == pht_waddr ? pht_5_34 : _GEN_3617; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3619 = 3'h5 == pht_windex & 6'h23 == pht_waddr ? pht_5_35 : _GEN_3618; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3620 = 3'h5 == pht_windex & 6'h24 == pht_waddr ? pht_5_36 : _GEN_3619; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3621 = 3'h5 == pht_windex & 6'h25 == pht_waddr ? pht_5_37 : _GEN_3620; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3622 = 3'h5 == pht_windex & 6'h26 == pht_waddr ? pht_5_38 : _GEN_3621; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3623 = 3'h5 == pht_windex & 6'h27 == pht_waddr ? pht_5_39 : _GEN_3622; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3624 = 3'h5 == pht_windex & 6'h28 == pht_waddr ? pht_5_40 : _GEN_3623; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3625 = 3'h5 == pht_windex & 6'h29 == pht_waddr ? pht_5_41 : _GEN_3624; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3626 = 3'h5 == pht_windex & 6'h2a == pht_waddr ? pht_5_42 : _GEN_3625; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3627 = 3'h5 == pht_windex & 6'h2b == pht_waddr ? pht_5_43 : _GEN_3626; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3628 = 3'h5 == pht_windex & 6'h2c == pht_waddr ? pht_5_44 : _GEN_3627; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3629 = 3'h5 == pht_windex & 6'h2d == pht_waddr ? pht_5_45 : _GEN_3628; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3630 = 3'h5 == pht_windex & 6'h2e == pht_waddr ? pht_5_46 : _GEN_3629; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3631 = 3'h5 == pht_windex & 6'h2f == pht_waddr ? pht_5_47 : _GEN_3630; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3632 = 3'h5 == pht_windex & 6'h30 == pht_waddr ? pht_5_48 : _GEN_3631; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3633 = 3'h5 == pht_windex & 6'h31 == pht_waddr ? pht_5_49 : _GEN_3632; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3634 = 3'h5 == pht_windex & 6'h32 == pht_waddr ? pht_5_50 : _GEN_3633; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3635 = 3'h5 == pht_windex & 6'h33 == pht_waddr ? pht_5_51 : _GEN_3634; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3636 = 3'h5 == pht_windex & 6'h34 == pht_waddr ? pht_5_52 : _GEN_3635; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3637 = 3'h5 == pht_windex & 6'h35 == pht_waddr ? pht_5_53 : _GEN_3636; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3638 = 3'h5 == pht_windex & 6'h36 == pht_waddr ? pht_5_54 : _GEN_3637; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3639 = 3'h5 == pht_windex & 6'h37 == pht_waddr ? pht_5_55 : _GEN_3638; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3640 = 3'h5 == pht_windex & 6'h38 == pht_waddr ? pht_5_56 : _GEN_3639; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3641 = 3'h5 == pht_windex & 6'h39 == pht_waddr ? pht_5_57 : _GEN_3640; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3642 = 3'h5 == pht_windex & 6'h3a == pht_waddr ? pht_5_58 : _GEN_3641; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3643 = 3'h5 == pht_windex & 6'h3b == pht_waddr ? pht_5_59 : _GEN_3642; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3644 = 3'h5 == pht_windex & 6'h3c == pht_waddr ? pht_5_60 : _GEN_3643; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3645 = 3'h5 == pht_windex & 6'h3d == pht_waddr ? pht_5_61 : _GEN_3644; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3646 = 3'h5 == pht_windex & 6'h3e == pht_waddr ? pht_5_62 : _GEN_3645; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3647 = 3'h5 == pht_windex & 6'h3f == pht_waddr ? pht_5_63 : _GEN_3646; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3648 = 3'h5 == pht_windex & 7'h40 == _GEN_14784 ? pht_5_64 : _GEN_3647; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3649 = 3'h5 == pht_windex & 7'h41 == _GEN_14784 ? pht_5_65 : _GEN_3648; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3650 = 3'h5 == pht_windex & 7'h42 == _GEN_14784 ? pht_5_66 : _GEN_3649; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3651 = 3'h5 == pht_windex & 7'h43 == _GEN_14784 ? pht_5_67 : _GEN_3650; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3652 = 3'h5 == pht_windex & 7'h44 == _GEN_14784 ? pht_5_68 : _GEN_3651; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3653 = 3'h5 == pht_windex & 7'h45 == _GEN_14784 ? pht_5_69 : _GEN_3652; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3654 = 3'h5 == pht_windex & 7'h46 == _GEN_14784 ? pht_5_70 : _GEN_3653; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3655 = 3'h5 == pht_windex & 7'h47 == _GEN_14784 ? pht_5_71 : _GEN_3654; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3656 = 3'h5 == pht_windex & 7'h48 == _GEN_14784 ? pht_5_72 : _GEN_3655; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3657 = 3'h5 == pht_windex & 7'h49 == _GEN_14784 ? pht_5_73 : _GEN_3656; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3658 = 3'h5 == pht_windex & 7'h4a == _GEN_14784 ? pht_5_74 : _GEN_3657; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3659 = 3'h5 == pht_windex & 7'h4b == _GEN_14784 ? pht_5_75 : _GEN_3658; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3660 = 3'h5 == pht_windex & 7'h4c == _GEN_14784 ? pht_5_76 : _GEN_3659; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3661 = 3'h5 == pht_windex & 7'h4d == _GEN_14784 ? pht_5_77 : _GEN_3660; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3662 = 3'h5 == pht_windex & 7'h4e == _GEN_14784 ? pht_5_78 : _GEN_3661; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3663 = 3'h5 == pht_windex & 7'h4f == _GEN_14784 ? pht_5_79 : _GEN_3662; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3664 = 3'h5 == pht_windex & 7'h50 == _GEN_14784 ? pht_5_80 : _GEN_3663; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3665 = 3'h5 == pht_windex & 7'h51 == _GEN_14784 ? pht_5_81 : _GEN_3664; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3666 = 3'h5 == pht_windex & 7'h52 == _GEN_14784 ? pht_5_82 : _GEN_3665; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3667 = 3'h5 == pht_windex & 7'h53 == _GEN_14784 ? pht_5_83 : _GEN_3666; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3668 = 3'h5 == pht_windex & 7'h54 == _GEN_14784 ? pht_5_84 : _GEN_3667; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3669 = 3'h5 == pht_windex & 7'h55 == _GEN_14784 ? pht_5_85 : _GEN_3668; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3670 = 3'h5 == pht_windex & 7'h56 == _GEN_14784 ? pht_5_86 : _GEN_3669; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3671 = 3'h5 == pht_windex & 7'h57 == _GEN_14784 ? pht_5_87 : _GEN_3670; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3672 = 3'h5 == pht_windex & 7'h58 == _GEN_14784 ? pht_5_88 : _GEN_3671; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3673 = 3'h5 == pht_windex & 7'h59 == _GEN_14784 ? pht_5_89 : _GEN_3672; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3674 = 3'h5 == pht_windex & 7'h5a == _GEN_14784 ? pht_5_90 : _GEN_3673; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3675 = 3'h5 == pht_windex & 7'h5b == _GEN_14784 ? pht_5_91 : _GEN_3674; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3676 = 3'h5 == pht_windex & 7'h5c == _GEN_14784 ? pht_5_92 : _GEN_3675; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3677 = 3'h5 == pht_windex & 7'h5d == _GEN_14784 ? pht_5_93 : _GEN_3676; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3678 = 3'h5 == pht_windex & 7'h5e == _GEN_14784 ? pht_5_94 : _GEN_3677; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3679 = 3'h5 == pht_windex & 7'h5f == _GEN_14784 ? pht_5_95 : _GEN_3678; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3680 = 3'h5 == pht_windex & 7'h60 == _GEN_14784 ? pht_5_96 : _GEN_3679; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3681 = 3'h5 == pht_windex & 7'h61 == _GEN_14784 ? pht_5_97 : _GEN_3680; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3682 = 3'h5 == pht_windex & 7'h62 == _GEN_14784 ? pht_5_98 : _GEN_3681; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3683 = 3'h5 == pht_windex & 7'h63 == _GEN_14784 ? pht_5_99 : _GEN_3682; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3684 = 3'h5 == pht_windex & 7'h64 == _GEN_14784 ? pht_5_100 : _GEN_3683; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3685 = 3'h5 == pht_windex & 7'h65 == _GEN_14784 ? pht_5_101 : _GEN_3684; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3686 = 3'h5 == pht_windex & 7'h66 == _GEN_14784 ? pht_5_102 : _GEN_3685; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3687 = 3'h5 == pht_windex & 7'h67 == _GEN_14784 ? pht_5_103 : _GEN_3686; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3688 = 3'h5 == pht_windex & 7'h68 == _GEN_14784 ? pht_5_104 : _GEN_3687; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3689 = 3'h5 == pht_windex & 7'h69 == _GEN_14784 ? pht_5_105 : _GEN_3688; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3690 = 3'h5 == pht_windex & 7'h6a == _GEN_14784 ? pht_5_106 : _GEN_3689; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3691 = 3'h5 == pht_windex & 7'h6b == _GEN_14784 ? pht_5_107 : _GEN_3690; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3692 = 3'h5 == pht_windex & 7'h6c == _GEN_14784 ? pht_5_108 : _GEN_3691; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3693 = 3'h5 == pht_windex & 7'h6d == _GEN_14784 ? pht_5_109 : _GEN_3692; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3694 = 3'h5 == pht_windex & 7'h6e == _GEN_14784 ? pht_5_110 : _GEN_3693; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3695 = 3'h5 == pht_windex & 7'h6f == _GEN_14784 ? pht_5_111 : _GEN_3694; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3696 = 3'h5 == pht_windex & 7'h70 == _GEN_14784 ? pht_5_112 : _GEN_3695; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3697 = 3'h5 == pht_windex & 7'h71 == _GEN_14784 ? pht_5_113 : _GEN_3696; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3698 = 3'h5 == pht_windex & 7'h72 == _GEN_14784 ? pht_5_114 : _GEN_3697; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3699 = 3'h5 == pht_windex & 7'h73 == _GEN_14784 ? pht_5_115 : _GEN_3698; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3700 = 3'h5 == pht_windex & 7'h74 == _GEN_14784 ? pht_5_116 : _GEN_3699; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3701 = 3'h5 == pht_windex & 7'h75 == _GEN_14784 ? pht_5_117 : _GEN_3700; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3702 = 3'h5 == pht_windex & 7'h76 == _GEN_14784 ? pht_5_118 : _GEN_3701; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3703 = 3'h5 == pht_windex & 7'h77 == _GEN_14784 ? pht_5_119 : _GEN_3702; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3704 = 3'h5 == pht_windex & 7'h78 == _GEN_14784 ? pht_5_120 : _GEN_3703; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3705 = 3'h5 == pht_windex & 7'h79 == _GEN_14784 ? pht_5_121 : _GEN_3704; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3706 = 3'h5 == pht_windex & 7'h7a == _GEN_14784 ? pht_5_122 : _GEN_3705; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3707 = 3'h5 == pht_windex & 7'h7b == _GEN_14784 ? pht_5_123 : _GEN_3706; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3708 = 3'h5 == pht_windex & 7'h7c == _GEN_14784 ? pht_5_124 : _GEN_3707; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3709 = 3'h5 == pht_windex & 7'h7d == _GEN_14784 ? pht_5_125 : _GEN_3708; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3710 = 3'h5 == pht_windex & 7'h7e == _GEN_14784 ? pht_5_126 : _GEN_3709; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3711 = 3'h5 == pht_windex & 7'h7f == _GEN_14784 ? pht_5_127 : _GEN_3710; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3712 = 3'h5 == pht_windex & 8'h80 == _GEN_14976 ? pht_5_128 : _GEN_3711; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3713 = 3'h5 == pht_windex & 8'h81 == _GEN_14976 ? pht_5_129 : _GEN_3712; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3714 = 3'h5 == pht_windex & 8'h82 == _GEN_14976 ? pht_5_130 : _GEN_3713; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3715 = 3'h5 == pht_windex & 8'h83 == _GEN_14976 ? pht_5_131 : _GEN_3714; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3716 = 3'h5 == pht_windex & 8'h84 == _GEN_14976 ? pht_5_132 : _GEN_3715; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3717 = 3'h5 == pht_windex & 8'h85 == _GEN_14976 ? pht_5_133 : _GEN_3716; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3718 = 3'h5 == pht_windex & 8'h86 == _GEN_14976 ? pht_5_134 : _GEN_3717; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3719 = 3'h5 == pht_windex & 8'h87 == _GEN_14976 ? pht_5_135 : _GEN_3718; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3720 = 3'h5 == pht_windex & 8'h88 == _GEN_14976 ? pht_5_136 : _GEN_3719; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3721 = 3'h5 == pht_windex & 8'h89 == _GEN_14976 ? pht_5_137 : _GEN_3720; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3722 = 3'h5 == pht_windex & 8'h8a == _GEN_14976 ? pht_5_138 : _GEN_3721; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3723 = 3'h5 == pht_windex & 8'h8b == _GEN_14976 ? pht_5_139 : _GEN_3722; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3724 = 3'h5 == pht_windex & 8'h8c == _GEN_14976 ? pht_5_140 : _GEN_3723; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3725 = 3'h5 == pht_windex & 8'h8d == _GEN_14976 ? pht_5_141 : _GEN_3724; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3726 = 3'h5 == pht_windex & 8'h8e == _GEN_14976 ? pht_5_142 : _GEN_3725; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3727 = 3'h5 == pht_windex & 8'h8f == _GEN_14976 ? pht_5_143 : _GEN_3726; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3728 = 3'h5 == pht_windex & 8'h90 == _GEN_14976 ? pht_5_144 : _GEN_3727; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3729 = 3'h5 == pht_windex & 8'h91 == _GEN_14976 ? pht_5_145 : _GEN_3728; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3730 = 3'h5 == pht_windex & 8'h92 == _GEN_14976 ? pht_5_146 : _GEN_3729; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3731 = 3'h5 == pht_windex & 8'h93 == _GEN_14976 ? pht_5_147 : _GEN_3730; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3732 = 3'h5 == pht_windex & 8'h94 == _GEN_14976 ? pht_5_148 : _GEN_3731; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3733 = 3'h5 == pht_windex & 8'h95 == _GEN_14976 ? pht_5_149 : _GEN_3732; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3734 = 3'h5 == pht_windex & 8'h96 == _GEN_14976 ? pht_5_150 : _GEN_3733; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3735 = 3'h5 == pht_windex & 8'h97 == _GEN_14976 ? pht_5_151 : _GEN_3734; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3736 = 3'h5 == pht_windex & 8'h98 == _GEN_14976 ? pht_5_152 : _GEN_3735; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3737 = 3'h5 == pht_windex & 8'h99 == _GEN_14976 ? pht_5_153 : _GEN_3736; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3738 = 3'h5 == pht_windex & 8'h9a == _GEN_14976 ? pht_5_154 : _GEN_3737; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3739 = 3'h5 == pht_windex & 8'h9b == _GEN_14976 ? pht_5_155 : _GEN_3738; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3740 = 3'h5 == pht_windex & 8'h9c == _GEN_14976 ? pht_5_156 : _GEN_3739; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3741 = 3'h5 == pht_windex & 8'h9d == _GEN_14976 ? pht_5_157 : _GEN_3740; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3742 = 3'h5 == pht_windex & 8'h9e == _GEN_14976 ? pht_5_158 : _GEN_3741; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3743 = 3'h5 == pht_windex & 8'h9f == _GEN_14976 ? pht_5_159 : _GEN_3742; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3744 = 3'h5 == pht_windex & 8'ha0 == _GEN_14976 ? pht_5_160 : _GEN_3743; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3745 = 3'h5 == pht_windex & 8'ha1 == _GEN_14976 ? pht_5_161 : _GEN_3744; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3746 = 3'h5 == pht_windex & 8'ha2 == _GEN_14976 ? pht_5_162 : _GEN_3745; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3747 = 3'h5 == pht_windex & 8'ha3 == _GEN_14976 ? pht_5_163 : _GEN_3746; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3748 = 3'h5 == pht_windex & 8'ha4 == _GEN_14976 ? pht_5_164 : _GEN_3747; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3749 = 3'h5 == pht_windex & 8'ha5 == _GEN_14976 ? pht_5_165 : _GEN_3748; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3750 = 3'h5 == pht_windex & 8'ha6 == _GEN_14976 ? pht_5_166 : _GEN_3749; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3751 = 3'h5 == pht_windex & 8'ha7 == _GEN_14976 ? pht_5_167 : _GEN_3750; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3752 = 3'h5 == pht_windex & 8'ha8 == _GEN_14976 ? pht_5_168 : _GEN_3751; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3753 = 3'h5 == pht_windex & 8'ha9 == _GEN_14976 ? pht_5_169 : _GEN_3752; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3754 = 3'h5 == pht_windex & 8'haa == _GEN_14976 ? pht_5_170 : _GEN_3753; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3755 = 3'h5 == pht_windex & 8'hab == _GEN_14976 ? pht_5_171 : _GEN_3754; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3756 = 3'h5 == pht_windex & 8'hac == _GEN_14976 ? pht_5_172 : _GEN_3755; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3757 = 3'h5 == pht_windex & 8'had == _GEN_14976 ? pht_5_173 : _GEN_3756; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3758 = 3'h5 == pht_windex & 8'hae == _GEN_14976 ? pht_5_174 : _GEN_3757; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3759 = 3'h5 == pht_windex & 8'haf == _GEN_14976 ? pht_5_175 : _GEN_3758; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3760 = 3'h5 == pht_windex & 8'hb0 == _GEN_14976 ? pht_5_176 : _GEN_3759; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3761 = 3'h5 == pht_windex & 8'hb1 == _GEN_14976 ? pht_5_177 : _GEN_3760; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3762 = 3'h5 == pht_windex & 8'hb2 == _GEN_14976 ? pht_5_178 : _GEN_3761; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3763 = 3'h5 == pht_windex & 8'hb3 == _GEN_14976 ? pht_5_179 : _GEN_3762; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3764 = 3'h5 == pht_windex & 8'hb4 == _GEN_14976 ? pht_5_180 : _GEN_3763; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3765 = 3'h5 == pht_windex & 8'hb5 == _GEN_14976 ? pht_5_181 : _GEN_3764; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3766 = 3'h5 == pht_windex & 8'hb6 == _GEN_14976 ? pht_5_182 : _GEN_3765; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3767 = 3'h5 == pht_windex & 8'hb7 == _GEN_14976 ? pht_5_183 : _GEN_3766; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3768 = 3'h5 == pht_windex & 8'hb8 == _GEN_14976 ? pht_5_184 : _GEN_3767; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3769 = 3'h5 == pht_windex & 8'hb9 == _GEN_14976 ? pht_5_185 : _GEN_3768; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3770 = 3'h5 == pht_windex & 8'hba == _GEN_14976 ? pht_5_186 : _GEN_3769; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3771 = 3'h5 == pht_windex & 8'hbb == _GEN_14976 ? pht_5_187 : _GEN_3770; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3772 = 3'h5 == pht_windex & 8'hbc == _GEN_14976 ? pht_5_188 : _GEN_3771; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3773 = 3'h5 == pht_windex & 8'hbd == _GEN_14976 ? pht_5_189 : _GEN_3772; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3774 = 3'h5 == pht_windex & 8'hbe == _GEN_14976 ? pht_5_190 : _GEN_3773; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3775 = 3'h5 == pht_windex & 8'hbf == _GEN_14976 ? pht_5_191 : _GEN_3774; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3776 = 3'h5 == pht_windex & 8'hc0 == _GEN_14976 ? pht_5_192 : _GEN_3775; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3777 = 3'h5 == pht_windex & 8'hc1 == _GEN_14976 ? pht_5_193 : _GEN_3776; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3778 = 3'h5 == pht_windex & 8'hc2 == _GEN_14976 ? pht_5_194 : _GEN_3777; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3779 = 3'h5 == pht_windex & 8'hc3 == _GEN_14976 ? pht_5_195 : _GEN_3778; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3780 = 3'h5 == pht_windex & 8'hc4 == _GEN_14976 ? pht_5_196 : _GEN_3779; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3781 = 3'h5 == pht_windex & 8'hc5 == _GEN_14976 ? pht_5_197 : _GEN_3780; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3782 = 3'h5 == pht_windex & 8'hc6 == _GEN_14976 ? pht_5_198 : _GEN_3781; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3783 = 3'h5 == pht_windex & 8'hc7 == _GEN_14976 ? pht_5_199 : _GEN_3782; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3784 = 3'h5 == pht_windex & 8'hc8 == _GEN_14976 ? pht_5_200 : _GEN_3783; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3785 = 3'h5 == pht_windex & 8'hc9 == _GEN_14976 ? pht_5_201 : _GEN_3784; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3786 = 3'h5 == pht_windex & 8'hca == _GEN_14976 ? pht_5_202 : _GEN_3785; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3787 = 3'h5 == pht_windex & 8'hcb == _GEN_14976 ? pht_5_203 : _GEN_3786; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3788 = 3'h5 == pht_windex & 8'hcc == _GEN_14976 ? pht_5_204 : _GEN_3787; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3789 = 3'h5 == pht_windex & 8'hcd == _GEN_14976 ? pht_5_205 : _GEN_3788; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3790 = 3'h5 == pht_windex & 8'hce == _GEN_14976 ? pht_5_206 : _GEN_3789; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3791 = 3'h5 == pht_windex & 8'hcf == _GEN_14976 ? pht_5_207 : _GEN_3790; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3792 = 3'h5 == pht_windex & 8'hd0 == _GEN_14976 ? pht_5_208 : _GEN_3791; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3793 = 3'h5 == pht_windex & 8'hd1 == _GEN_14976 ? pht_5_209 : _GEN_3792; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3794 = 3'h5 == pht_windex & 8'hd2 == _GEN_14976 ? pht_5_210 : _GEN_3793; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3795 = 3'h5 == pht_windex & 8'hd3 == _GEN_14976 ? pht_5_211 : _GEN_3794; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3796 = 3'h5 == pht_windex & 8'hd4 == _GEN_14976 ? pht_5_212 : _GEN_3795; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3797 = 3'h5 == pht_windex & 8'hd5 == _GEN_14976 ? pht_5_213 : _GEN_3796; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3798 = 3'h5 == pht_windex & 8'hd6 == _GEN_14976 ? pht_5_214 : _GEN_3797; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3799 = 3'h5 == pht_windex & 8'hd7 == _GEN_14976 ? pht_5_215 : _GEN_3798; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3800 = 3'h5 == pht_windex & 8'hd8 == _GEN_14976 ? pht_5_216 : _GEN_3799; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3801 = 3'h5 == pht_windex & 8'hd9 == _GEN_14976 ? pht_5_217 : _GEN_3800; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3802 = 3'h5 == pht_windex & 8'hda == _GEN_14976 ? pht_5_218 : _GEN_3801; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3803 = 3'h5 == pht_windex & 8'hdb == _GEN_14976 ? pht_5_219 : _GEN_3802; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3804 = 3'h5 == pht_windex & 8'hdc == _GEN_14976 ? pht_5_220 : _GEN_3803; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3805 = 3'h5 == pht_windex & 8'hdd == _GEN_14976 ? pht_5_221 : _GEN_3804; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3806 = 3'h5 == pht_windex & 8'hde == _GEN_14976 ? pht_5_222 : _GEN_3805; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3807 = 3'h5 == pht_windex & 8'hdf == _GEN_14976 ? pht_5_223 : _GEN_3806; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3808 = 3'h5 == pht_windex & 8'he0 == _GEN_14976 ? pht_5_224 : _GEN_3807; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3809 = 3'h5 == pht_windex & 8'he1 == _GEN_14976 ? pht_5_225 : _GEN_3808; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3810 = 3'h5 == pht_windex & 8'he2 == _GEN_14976 ? pht_5_226 : _GEN_3809; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3811 = 3'h5 == pht_windex & 8'he3 == _GEN_14976 ? pht_5_227 : _GEN_3810; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3812 = 3'h5 == pht_windex & 8'he4 == _GEN_14976 ? pht_5_228 : _GEN_3811; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3813 = 3'h5 == pht_windex & 8'he5 == _GEN_14976 ? pht_5_229 : _GEN_3812; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3814 = 3'h5 == pht_windex & 8'he6 == _GEN_14976 ? pht_5_230 : _GEN_3813; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3815 = 3'h5 == pht_windex & 8'he7 == _GEN_14976 ? pht_5_231 : _GEN_3814; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3816 = 3'h5 == pht_windex & 8'he8 == _GEN_14976 ? pht_5_232 : _GEN_3815; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3817 = 3'h5 == pht_windex & 8'he9 == _GEN_14976 ? pht_5_233 : _GEN_3816; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3818 = 3'h5 == pht_windex & 8'hea == _GEN_14976 ? pht_5_234 : _GEN_3817; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3819 = 3'h5 == pht_windex & 8'heb == _GEN_14976 ? pht_5_235 : _GEN_3818; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3820 = 3'h5 == pht_windex & 8'hec == _GEN_14976 ? pht_5_236 : _GEN_3819; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3821 = 3'h5 == pht_windex & 8'hed == _GEN_14976 ? pht_5_237 : _GEN_3820; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3822 = 3'h5 == pht_windex & 8'hee == _GEN_14976 ? pht_5_238 : _GEN_3821; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3823 = 3'h5 == pht_windex & 8'hef == _GEN_14976 ? pht_5_239 : _GEN_3822; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3824 = 3'h5 == pht_windex & 8'hf0 == _GEN_14976 ? pht_5_240 : _GEN_3823; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3825 = 3'h5 == pht_windex & 8'hf1 == _GEN_14976 ? pht_5_241 : _GEN_3824; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3826 = 3'h5 == pht_windex & 8'hf2 == _GEN_14976 ? pht_5_242 : _GEN_3825; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3827 = 3'h5 == pht_windex & 8'hf3 == _GEN_14976 ? pht_5_243 : _GEN_3826; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3828 = 3'h5 == pht_windex & 8'hf4 == _GEN_14976 ? pht_5_244 : _GEN_3827; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3829 = 3'h5 == pht_windex & 8'hf5 == _GEN_14976 ? pht_5_245 : _GEN_3828; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3830 = 3'h5 == pht_windex & 8'hf6 == _GEN_14976 ? pht_5_246 : _GEN_3829; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3831 = 3'h5 == pht_windex & 8'hf7 == _GEN_14976 ? pht_5_247 : _GEN_3830; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3832 = 3'h5 == pht_windex & 8'hf8 == _GEN_14976 ? pht_5_248 : _GEN_3831; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3833 = 3'h5 == pht_windex & 8'hf9 == _GEN_14976 ? pht_5_249 : _GEN_3832; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3834 = 3'h5 == pht_windex & 8'hfa == _GEN_14976 ? pht_5_250 : _GEN_3833; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3835 = 3'h5 == pht_windex & 8'hfb == _GEN_14976 ? pht_5_251 : _GEN_3834; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3836 = 3'h5 == pht_windex & 8'hfc == _GEN_14976 ? pht_5_252 : _GEN_3835; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3837 = 3'h5 == pht_windex & 8'hfd == _GEN_14976 ? pht_5_253 : _GEN_3836; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3838 = 3'h5 == pht_windex & 8'hfe == _GEN_14976 ? pht_5_254 : _GEN_3837; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3839 = 3'h5 == pht_windex & 8'hff == _GEN_14976 ? pht_5_255 : _GEN_3838; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_18880 = 3'h6 == pht_windex; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3840 = 3'h6 == pht_windex & 6'h0 == pht_waddr ? pht_6_0 : _GEN_3839; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3841 = 3'h6 == pht_windex & 6'h1 == pht_waddr ? pht_6_1 : _GEN_3840; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3842 = 3'h6 == pht_windex & 6'h2 == pht_waddr ? pht_6_2 : _GEN_3841; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3843 = 3'h6 == pht_windex & 6'h3 == pht_waddr ? pht_6_3 : _GEN_3842; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3844 = 3'h6 == pht_windex & 6'h4 == pht_waddr ? pht_6_4 : _GEN_3843; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3845 = 3'h6 == pht_windex & 6'h5 == pht_waddr ? pht_6_5 : _GEN_3844; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3846 = 3'h6 == pht_windex & 6'h6 == pht_waddr ? pht_6_6 : _GEN_3845; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3847 = 3'h6 == pht_windex & 6'h7 == pht_waddr ? pht_6_7 : _GEN_3846; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3848 = 3'h6 == pht_windex & 6'h8 == pht_waddr ? pht_6_8 : _GEN_3847; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3849 = 3'h6 == pht_windex & 6'h9 == pht_waddr ? pht_6_9 : _GEN_3848; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3850 = 3'h6 == pht_windex & 6'ha == pht_waddr ? pht_6_10 : _GEN_3849; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3851 = 3'h6 == pht_windex & 6'hb == pht_waddr ? pht_6_11 : _GEN_3850; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3852 = 3'h6 == pht_windex & 6'hc == pht_waddr ? pht_6_12 : _GEN_3851; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3853 = 3'h6 == pht_windex & 6'hd == pht_waddr ? pht_6_13 : _GEN_3852; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3854 = 3'h6 == pht_windex & 6'he == pht_waddr ? pht_6_14 : _GEN_3853; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3855 = 3'h6 == pht_windex & 6'hf == pht_waddr ? pht_6_15 : _GEN_3854; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3856 = 3'h6 == pht_windex & 6'h10 == pht_waddr ? pht_6_16 : _GEN_3855; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3857 = 3'h6 == pht_windex & 6'h11 == pht_waddr ? pht_6_17 : _GEN_3856; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3858 = 3'h6 == pht_windex & 6'h12 == pht_waddr ? pht_6_18 : _GEN_3857; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3859 = 3'h6 == pht_windex & 6'h13 == pht_waddr ? pht_6_19 : _GEN_3858; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3860 = 3'h6 == pht_windex & 6'h14 == pht_waddr ? pht_6_20 : _GEN_3859; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3861 = 3'h6 == pht_windex & 6'h15 == pht_waddr ? pht_6_21 : _GEN_3860; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3862 = 3'h6 == pht_windex & 6'h16 == pht_waddr ? pht_6_22 : _GEN_3861; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3863 = 3'h6 == pht_windex & 6'h17 == pht_waddr ? pht_6_23 : _GEN_3862; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3864 = 3'h6 == pht_windex & 6'h18 == pht_waddr ? pht_6_24 : _GEN_3863; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3865 = 3'h6 == pht_windex & 6'h19 == pht_waddr ? pht_6_25 : _GEN_3864; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3866 = 3'h6 == pht_windex & 6'h1a == pht_waddr ? pht_6_26 : _GEN_3865; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3867 = 3'h6 == pht_windex & 6'h1b == pht_waddr ? pht_6_27 : _GEN_3866; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3868 = 3'h6 == pht_windex & 6'h1c == pht_waddr ? pht_6_28 : _GEN_3867; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3869 = 3'h6 == pht_windex & 6'h1d == pht_waddr ? pht_6_29 : _GEN_3868; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3870 = 3'h6 == pht_windex & 6'h1e == pht_waddr ? pht_6_30 : _GEN_3869; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3871 = 3'h6 == pht_windex & 6'h1f == pht_waddr ? pht_6_31 : _GEN_3870; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3872 = 3'h6 == pht_windex & 6'h20 == pht_waddr ? pht_6_32 : _GEN_3871; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3873 = 3'h6 == pht_windex & 6'h21 == pht_waddr ? pht_6_33 : _GEN_3872; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3874 = 3'h6 == pht_windex & 6'h22 == pht_waddr ? pht_6_34 : _GEN_3873; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3875 = 3'h6 == pht_windex & 6'h23 == pht_waddr ? pht_6_35 : _GEN_3874; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3876 = 3'h6 == pht_windex & 6'h24 == pht_waddr ? pht_6_36 : _GEN_3875; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3877 = 3'h6 == pht_windex & 6'h25 == pht_waddr ? pht_6_37 : _GEN_3876; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3878 = 3'h6 == pht_windex & 6'h26 == pht_waddr ? pht_6_38 : _GEN_3877; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3879 = 3'h6 == pht_windex & 6'h27 == pht_waddr ? pht_6_39 : _GEN_3878; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3880 = 3'h6 == pht_windex & 6'h28 == pht_waddr ? pht_6_40 : _GEN_3879; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3881 = 3'h6 == pht_windex & 6'h29 == pht_waddr ? pht_6_41 : _GEN_3880; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3882 = 3'h6 == pht_windex & 6'h2a == pht_waddr ? pht_6_42 : _GEN_3881; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3883 = 3'h6 == pht_windex & 6'h2b == pht_waddr ? pht_6_43 : _GEN_3882; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3884 = 3'h6 == pht_windex & 6'h2c == pht_waddr ? pht_6_44 : _GEN_3883; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3885 = 3'h6 == pht_windex & 6'h2d == pht_waddr ? pht_6_45 : _GEN_3884; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3886 = 3'h6 == pht_windex & 6'h2e == pht_waddr ? pht_6_46 : _GEN_3885; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3887 = 3'h6 == pht_windex & 6'h2f == pht_waddr ? pht_6_47 : _GEN_3886; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3888 = 3'h6 == pht_windex & 6'h30 == pht_waddr ? pht_6_48 : _GEN_3887; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3889 = 3'h6 == pht_windex & 6'h31 == pht_waddr ? pht_6_49 : _GEN_3888; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3890 = 3'h6 == pht_windex & 6'h32 == pht_waddr ? pht_6_50 : _GEN_3889; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3891 = 3'h6 == pht_windex & 6'h33 == pht_waddr ? pht_6_51 : _GEN_3890; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3892 = 3'h6 == pht_windex & 6'h34 == pht_waddr ? pht_6_52 : _GEN_3891; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3893 = 3'h6 == pht_windex & 6'h35 == pht_waddr ? pht_6_53 : _GEN_3892; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3894 = 3'h6 == pht_windex & 6'h36 == pht_waddr ? pht_6_54 : _GEN_3893; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3895 = 3'h6 == pht_windex & 6'h37 == pht_waddr ? pht_6_55 : _GEN_3894; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3896 = 3'h6 == pht_windex & 6'h38 == pht_waddr ? pht_6_56 : _GEN_3895; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3897 = 3'h6 == pht_windex & 6'h39 == pht_waddr ? pht_6_57 : _GEN_3896; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3898 = 3'h6 == pht_windex & 6'h3a == pht_waddr ? pht_6_58 : _GEN_3897; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3899 = 3'h6 == pht_windex & 6'h3b == pht_waddr ? pht_6_59 : _GEN_3898; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3900 = 3'h6 == pht_windex & 6'h3c == pht_waddr ? pht_6_60 : _GEN_3899; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3901 = 3'h6 == pht_windex & 6'h3d == pht_waddr ? pht_6_61 : _GEN_3900; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3902 = 3'h6 == pht_windex & 6'h3e == pht_waddr ? pht_6_62 : _GEN_3901; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3903 = 3'h6 == pht_windex & 6'h3f == pht_waddr ? pht_6_63 : _GEN_3902; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3904 = 3'h6 == pht_windex & 7'h40 == _GEN_14784 ? pht_6_64 : _GEN_3903; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3905 = 3'h6 == pht_windex & 7'h41 == _GEN_14784 ? pht_6_65 : _GEN_3904; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3906 = 3'h6 == pht_windex & 7'h42 == _GEN_14784 ? pht_6_66 : _GEN_3905; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3907 = 3'h6 == pht_windex & 7'h43 == _GEN_14784 ? pht_6_67 : _GEN_3906; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3908 = 3'h6 == pht_windex & 7'h44 == _GEN_14784 ? pht_6_68 : _GEN_3907; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3909 = 3'h6 == pht_windex & 7'h45 == _GEN_14784 ? pht_6_69 : _GEN_3908; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3910 = 3'h6 == pht_windex & 7'h46 == _GEN_14784 ? pht_6_70 : _GEN_3909; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3911 = 3'h6 == pht_windex & 7'h47 == _GEN_14784 ? pht_6_71 : _GEN_3910; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3912 = 3'h6 == pht_windex & 7'h48 == _GEN_14784 ? pht_6_72 : _GEN_3911; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3913 = 3'h6 == pht_windex & 7'h49 == _GEN_14784 ? pht_6_73 : _GEN_3912; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3914 = 3'h6 == pht_windex & 7'h4a == _GEN_14784 ? pht_6_74 : _GEN_3913; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3915 = 3'h6 == pht_windex & 7'h4b == _GEN_14784 ? pht_6_75 : _GEN_3914; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3916 = 3'h6 == pht_windex & 7'h4c == _GEN_14784 ? pht_6_76 : _GEN_3915; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3917 = 3'h6 == pht_windex & 7'h4d == _GEN_14784 ? pht_6_77 : _GEN_3916; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3918 = 3'h6 == pht_windex & 7'h4e == _GEN_14784 ? pht_6_78 : _GEN_3917; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3919 = 3'h6 == pht_windex & 7'h4f == _GEN_14784 ? pht_6_79 : _GEN_3918; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3920 = 3'h6 == pht_windex & 7'h50 == _GEN_14784 ? pht_6_80 : _GEN_3919; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3921 = 3'h6 == pht_windex & 7'h51 == _GEN_14784 ? pht_6_81 : _GEN_3920; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3922 = 3'h6 == pht_windex & 7'h52 == _GEN_14784 ? pht_6_82 : _GEN_3921; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3923 = 3'h6 == pht_windex & 7'h53 == _GEN_14784 ? pht_6_83 : _GEN_3922; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3924 = 3'h6 == pht_windex & 7'h54 == _GEN_14784 ? pht_6_84 : _GEN_3923; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3925 = 3'h6 == pht_windex & 7'h55 == _GEN_14784 ? pht_6_85 : _GEN_3924; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3926 = 3'h6 == pht_windex & 7'h56 == _GEN_14784 ? pht_6_86 : _GEN_3925; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3927 = 3'h6 == pht_windex & 7'h57 == _GEN_14784 ? pht_6_87 : _GEN_3926; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3928 = 3'h6 == pht_windex & 7'h58 == _GEN_14784 ? pht_6_88 : _GEN_3927; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3929 = 3'h6 == pht_windex & 7'h59 == _GEN_14784 ? pht_6_89 : _GEN_3928; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3930 = 3'h6 == pht_windex & 7'h5a == _GEN_14784 ? pht_6_90 : _GEN_3929; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3931 = 3'h6 == pht_windex & 7'h5b == _GEN_14784 ? pht_6_91 : _GEN_3930; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3932 = 3'h6 == pht_windex & 7'h5c == _GEN_14784 ? pht_6_92 : _GEN_3931; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3933 = 3'h6 == pht_windex & 7'h5d == _GEN_14784 ? pht_6_93 : _GEN_3932; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3934 = 3'h6 == pht_windex & 7'h5e == _GEN_14784 ? pht_6_94 : _GEN_3933; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3935 = 3'h6 == pht_windex & 7'h5f == _GEN_14784 ? pht_6_95 : _GEN_3934; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3936 = 3'h6 == pht_windex & 7'h60 == _GEN_14784 ? pht_6_96 : _GEN_3935; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3937 = 3'h6 == pht_windex & 7'h61 == _GEN_14784 ? pht_6_97 : _GEN_3936; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3938 = 3'h6 == pht_windex & 7'h62 == _GEN_14784 ? pht_6_98 : _GEN_3937; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3939 = 3'h6 == pht_windex & 7'h63 == _GEN_14784 ? pht_6_99 : _GEN_3938; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3940 = 3'h6 == pht_windex & 7'h64 == _GEN_14784 ? pht_6_100 : _GEN_3939; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3941 = 3'h6 == pht_windex & 7'h65 == _GEN_14784 ? pht_6_101 : _GEN_3940; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3942 = 3'h6 == pht_windex & 7'h66 == _GEN_14784 ? pht_6_102 : _GEN_3941; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3943 = 3'h6 == pht_windex & 7'h67 == _GEN_14784 ? pht_6_103 : _GEN_3942; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3944 = 3'h6 == pht_windex & 7'h68 == _GEN_14784 ? pht_6_104 : _GEN_3943; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3945 = 3'h6 == pht_windex & 7'h69 == _GEN_14784 ? pht_6_105 : _GEN_3944; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3946 = 3'h6 == pht_windex & 7'h6a == _GEN_14784 ? pht_6_106 : _GEN_3945; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3947 = 3'h6 == pht_windex & 7'h6b == _GEN_14784 ? pht_6_107 : _GEN_3946; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3948 = 3'h6 == pht_windex & 7'h6c == _GEN_14784 ? pht_6_108 : _GEN_3947; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3949 = 3'h6 == pht_windex & 7'h6d == _GEN_14784 ? pht_6_109 : _GEN_3948; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3950 = 3'h6 == pht_windex & 7'h6e == _GEN_14784 ? pht_6_110 : _GEN_3949; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3951 = 3'h6 == pht_windex & 7'h6f == _GEN_14784 ? pht_6_111 : _GEN_3950; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3952 = 3'h6 == pht_windex & 7'h70 == _GEN_14784 ? pht_6_112 : _GEN_3951; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3953 = 3'h6 == pht_windex & 7'h71 == _GEN_14784 ? pht_6_113 : _GEN_3952; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3954 = 3'h6 == pht_windex & 7'h72 == _GEN_14784 ? pht_6_114 : _GEN_3953; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3955 = 3'h6 == pht_windex & 7'h73 == _GEN_14784 ? pht_6_115 : _GEN_3954; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3956 = 3'h6 == pht_windex & 7'h74 == _GEN_14784 ? pht_6_116 : _GEN_3955; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3957 = 3'h6 == pht_windex & 7'h75 == _GEN_14784 ? pht_6_117 : _GEN_3956; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3958 = 3'h6 == pht_windex & 7'h76 == _GEN_14784 ? pht_6_118 : _GEN_3957; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3959 = 3'h6 == pht_windex & 7'h77 == _GEN_14784 ? pht_6_119 : _GEN_3958; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3960 = 3'h6 == pht_windex & 7'h78 == _GEN_14784 ? pht_6_120 : _GEN_3959; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3961 = 3'h6 == pht_windex & 7'h79 == _GEN_14784 ? pht_6_121 : _GEN_3960; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3962 = 3'h6 == pht_windex & 7'h7a == _GEN_14784 ? pht_6_122 : _GEN_3961; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3963 = 3'h6 == pht_windex & 7'h7b == _GEN_14784 ? pht_6_123 : _GEN_3962; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3964 = 3'h6 == pht_windex & 7'h7c == _GEN_14784 ? pht_6_124 : _GEN_3963; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3965 = 3'h6 == pht_windex & 7'h7d == _GEN_14784 ? pht_6_125 : _GEN_3964; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3966 = 3'h6 == pht_windex & 7'h7e == _GEN_14784 ? pht_6_126 : _GEN_3965; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3967 = 3'h6 == pht_windex & 7'h7f == _GEN_14784 ? pht_6_127 : _GEN_3966; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3968 = 3'h6 == pht_windex & 8'h80 == _GEN_14976 ? pht_6_128 : _GEN_3967; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3969 = 3'h6 == pht_windex & 8'h81 == _GEN_14976 ? pht_6_129 : _GEN_3968; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3970 = 3'h6 == pht_windex & 8'h82 == _GEN_14976 ? pht_6_130 : _GEN_3969; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3971 = 3'h6 == pht_windex & 8'h83 == _GEN_14976 ? pht_6_131 : _GEN_3970; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3972 = 3'h6 == pht_windex & 8'h84 == _GEN_14976 ? pht_6_132 : _GEN_3971; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3973 = 3'h6 == pht_windex & 8'h85 == _GEN_14976 ? pht_6_133 : _GEN_3972; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3974 = 3'h6 == pht_windex & 8'h86 == _GEN_14976 ? pht_6_134 : _GEN_3973; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3975 = 3'h6 == pht_windex & 8'h87 == _GEN_14976 ? pht_6_135 : _GEN_3974; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3976 = 3'h6 == pht_windex & 8'h88 == _GEN_14976 ? pht_6_136 : _GEN_3975; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3977 = 3'h6 == pht_windex & 8'h89 == _GEN_14976 ? pht_6_137 : _GEN_3976; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3978 = 3'h6 == pht_windex & 8'h8a == _GEN_14976 ? pht_6_138 : _GEN_3977; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3979 = 3'h6 == pht_windex & 8'h8b == _GEN_14976 ? pht_6_139 : _GEN_3978; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3980 = 3'h6 == pht_windex & 8'h8c == _GEN_14976 ? pht_6_140 : _GEN_3979; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3981 = 3'h6 == pht_windex & 8'h8d == _GEN_14976 ? pht_6_141 : _GEN_3980; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3982 = 3'h6 == pht_windex & 8'h8e == _GEN_14976 ? pht_6_142 : _GEN_3981; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3983 = 3'h6 == pht_windex & 8'h8f == _GEN_14976 ? pht_6_143 : _GEN_3982; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3984 = 3'h6 == pht_windex & 8'h90 == _GEN_14976 ? pht_6_144 : _GEN_3983; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3985 = 3'h6 == pht_windex & 8'h91 == _GEN_14976 ? pht_6_145 : _GEN_3984; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3986 = 3'h6 == pht_windex & 8'h92 == _GEN_14976 ? pht_6_146 : _GEN_3985; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3987 = 3'h6 == pht_windex & 8'h93 == _GEN_14976 ? pht_6_147 : _GEN_3986; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3988 = 3'h6 == pht_windex & 8'h94 == _GEN_14976 ? pht_6_148 : _GEN_3987; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3989 = 3'h6 == pht_windex & 8'h95 == _GEN_14976 ? pht_6_149 : _GEN_3988; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3990 = 3'h6 == pht_windex & 8'h96 == _GEN_14976 ? pht_6_150 : _GEN_3989; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3991 = 3'h6 == pht_windex & 8'h97 == _GEN_14976 ? pht_6_151 : _GEN_3990; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3992 = 3'h6 == pht_windex & 8'h98 == _GEN_14976 ? pht_6_152 : _GEN_3991; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3993 = 3'h6 == pht_windex & 8'h99 == _GEN_14976 ? pht_6_153 : _GEN_3992; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3994 = 3'h6 == pht_windex & 8'h9a == _GEN_14976 ? pht_6_154 : _GEN_3993; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3995 = 3'h6 == pht_windex & 8'h9b == _GEN_14976 ? pht_6_155 : _GEN_3994; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3996 = 3'h6 == pht_windex & 8'h9c == _GEN_14976 ? pht_6_156 : _GEN_3995; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3997 = 3'h6 == pht_windex & 8'h9d == _GEN_14976 ? pht_6_157 : _GEN_3996; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3998 = 3'h6 == pht_windex & 8'h9e == _GEN_14976 ? pht_6_158 : _GEN_3997; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_3999 = 3'h6 == pht_windex & 8'h9f == _GEN_14976 ? pht_6_159 : _GEN_3998; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4000 = 3'h6 == pht_windex & 8'ha0 == _GEN_14976 ? pht_6_160 : _GEN_3999; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4001 = 3'h6 == pht_windex & 8'ha1 == _GEN_14976 ? pht_6_161 : _GEN_4000; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4002 = 3'h6 == pht_windex & 8'ha2 == _GEN_14976 ? pht_6_162 : _GEN_4001; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4003 = 3'h6 == pht_windex & 8'ha3 == _GEN_14976 ? pht_6_163 : _GEN_4002; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4004 = 3'h6 == pht_windex & 8'ha4 == _GEN_14976 ? pht_6_164 : _GEN_4003; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4005 = 3'h6 == pht_windex & 8'ha5 == _GEN_14976 ? pht_6_165 : _GEN_4004; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4006 = 3'h6 == pht_windex & 8'ha6 == _GEN_14976 ? pht_6_166 : _GEN_4005; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4007 = 3'h6 == pht_windex & 8'ha7 == _GEN_14976 ? pht_6_167 : _GEN_4006; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4008 = 3'h6 == pht_windex & 8'ha8 == _GEN_14976 ? pht_6_168 : _GEN_4007; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4009 = 3'h6 == pht_windex & 8'ha9 == _GEN_14976 ? pht_6_169 : _GEN_4008; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4010 = 3'h6 == pht_windex & 8'haa == _GEN_14976 ? pht_6_170 : _GEN_4009; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4011 = 3'h6 == pht_windex & 8'hab == _GEN_14976 ? pht_6_171 : _GEN_4010; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4012 = 3'h6 == pht_windex & 8'hac == _GEN_14976 ? pht_6_172 : _GEN_4011; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4013 = 3'h6 == pht_windex & 8'had == _GEN_14976 ? pht_6_173 : _GEN_4012; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4014 = 3'h6 == pht_windex & 8'hae == _GEN_14976 ? pht_6_174 : _GEN_4013; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4015 = 3'h6 == pht_windex & 8'haf == _GEN_14976 ? pht_6_175 : _GEN_4014; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4016 = 3'h6 == pht_windex & 8'hb0 == _GEN_14976 ? pht_6_176 : _GEN_4015; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4017 = 3'h6 == pht_windex & 8'hb1 == _GEN_14976 ? pht_6_177 : _GEN_4016; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4018 = 3'h6 == pht_windex & 8'hb2 == _GEN_14976 ? pht_6_178 : _GEN_4017; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4019 = 3'h6 == pht_windex & 8'hb3 == _GEN_14976 ? pht_6_179 : _GEN_4018; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4020 = 3'h6 == pht_windex & 8'hb4 == _GEN_14976 ? pht_6_180 : _GEN_4019; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4021 = 3'h6 == pht_windex & 8'hb5 == _GEN_14976 ? pht_6_181 : _GEN_4020; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4022 = 3'h6 == pht_windex & 8'hb6 == _GEN_14976 ? pht_6_182 : _GEN_4021; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4023 = 3'h6 == pht_windex & 8'hb7 == _GEN_14976 ? pht_6_183 : _GEN_4022; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4024 = 3'h6 == pht_windex & 8'hb8 == _GEN_14976 ? pht_6_184 : _GEN_4023; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4025 = 3'h6 == pht_windex & 8'hb9 == _GEN_14976 ? pht_6_185 : _GEN_4024; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4026 = 3'h6 == pht_windex & 8'hba == _GEN_14976 ? pht_6_186 : _GEN_4025; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4027 = 3'h6 == pht_windex & 8'hbb == _GEN_14976 ? pht_6_187 : _GEN_4026; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4028 = 3'h6 == pht_windex & 8'hbc == _GEN_14976 ? pht_6_188 : _GEN_4027; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4029 = 3'h6 == pht_windex & 8'hbd == _GEN_14976 ? pht_6_189 : _GEN_4028; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4030 = 3'h6 == pht_windex & 8'hbe == _GEN_14976 ? pht_6_190 : _GEN_4029; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4031 = 3'h6 == pht_windex & 8'hbf == _GEN_14976 ? pht_6_191 : _GEN_4030; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4032 = 3'h6 == pht_windex & 8'hc0 == _GEN_14976 ? pht_6_192 : _GEN_4031; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4033 = 3'h6 == pht_windex & 8'hc1 == _GEN_14976 ? pht_6_193 : _GEN_4032; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4034 = 3'h6 == pht_windex & 8'hc2 == _GEN_14976 ? pht_6_194 : _GEN_4033; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4035 = 3'h6 == pht_windex & 8'hc3 == _GEN_14976 ? pht_6_195 : _GEN_4034; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4036 = 3'h6 == pht_windex & 8'hc4 == _GEN_14976 ? pht_6_196 : _GEN_4035; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4037 = 3'h6 == pht_windex & 8'hc5 == _GEN_14976 ? pht_6_197 : _GEN_4036; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4038 = 3'h6 == pht_windex & 8'hc6 == _GEN_14976 ? pht_6_198 : _GEN_4037; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4039 = 3'h6 == pht_windex & 8'hc7 == _GEN_14976 ? pht_6_199 : _GEN_4038; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4040 = 3'h6 == pht_windex & 8'hc8 == _GEN_14976 ? pht_6_200 : _GEN_4039; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4041 = 3'h6 == pht_windex & 8'hc9 == _GEN_14976 ? pht_6_201 : _GEN_4040; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4042 = 3'h6 == pht_windex & 8'hca == _GEN_14976 ? pht_6_202 : _GEN_4041; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4043 = 3'h6 == pht_windex & 8'hcb == _GEN_14976 ? pht_6_203 : _GEN_4042; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4044 = 3'h6 == pht_windex & 8'hcc == _GEN_14976 ? pht_6_204 : _GEN_4043; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4045 = 3'h6 == pht_windex & 8'hcd == _GEN_14976 ? pht_6_205 : _GEN_4044; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4046 = 3'h6 == pht_windex & 8'hce == _GEN_14976 ? pht_6_206 : _GEN_4045; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4047 = 3'h6 == pht_windex & 8'hcf == _GEN_14976 ? pht_6_207 : _GEN_4046; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4048 = 3'h6 == pht_windex & 8'hd0 == _GEN_14976 ? pht_6_208 : _GEN_4047; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4049 = 3'h6 == pht_windex & 8'hd1 == _GEN_14976 ? pht_6_209 : _GEN_4048; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4050 = 3'h6 == pht_windex & 8'hd2 == _GEN_14976 ? pht_6_210 : _GEN_4049; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4051 = 3'h6 == pht_windex & 8'hd3 == _GEN_14976 ? pht_6_211 : _GEN_4050; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4052 = 3'h6 == pht_windex & 8'hd4 == _GEN_14976 ? pht_6_212 : _GEN_4051; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4053 = 3'h6 == pht_windex & 8'hd5 == _GEN_14976 ? pht_6_213 : _GEN_4052; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4054 = 3'h6 == pht_windex & 8'hd6 == _GEN_14976 ? pht_6_214 : _GEN_4053; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4055 = 3'h6 == pht_windex & 8'hd7 == _GEN_14976 ? pht_6_215 : _GEN_4054; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4056 = 3'h6 == pht_windex & 8'hd8 == _GEN_14976 ? pht_6_216 : _GEN_4055; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4057 = 3'h6 == pht_windex & 8'hd9 == _GEN_14976 ? pht_6_217 : _GEN_4056; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4058 = 3'h6 == pht_windex & 8'hda == _GEN_14976 ? pht_6_218 : _GEN_4057; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4059 = 3'h6 == pht_windex & 8'hdb == _GEN_14976 ? pht_6_219 : _GEN_4058; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4060 = 3'h6 == pht_windex & 8'hdc == _GEN_14976 ? pht_6_220 : _GEN_4059; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4061 = 3'h6 == pht_windex & 8'hdd == _GEN_14976 ? pht_6_221 : _GEN_4060; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4062 = 3'h6 == pht_windex & 8'hde == _GEN_14976 ? pht_6_222 : _GEN_4061; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4063 = 3'h6 == pht_windex & 8'hdf == _GEN_14976 ? pht_6_223 : _GEN_4062; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4064 = 3'h6 == pht_windex & 8'he0 == _GEN_14976 ? pht_6_224 : _GEN_4063; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4065 = 3'h6 == pht_windex & 8'he1 == _GEN_14976 ? pht_6_225 : _GEN_4064; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4066 = 3'h6 == pht_windex & 8'he2 == _GEN_14976 ? pht_6_226 : _GEN_4065; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4067 = 3'h6 == pht_windex & 8'he3 == _GEN_14976 ? pht_6_227 : _GEN_4066; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4068 = 3'h6 == pht_windex & 8'he4 == _GEN_14976 ? pht_6_228 : _GEN_4067; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4069 = 3'h6 == pht_windex & 8'he5 == _GEN_14976 ? pht_6_229 : _GEN_4068; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4070 = 3'h6 == pht_windex & 8'he6 == _GEN_14976 ? pht_6_230 : _GEN_4069; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4071 = 3'h6 == pht_windex & 8'he7 == _GEN_14976 ? pht_6_231 : _GEN_4070; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4072 = 3'h6 == pht_windex & 8'he8 == _GEN_14976 ? pht_6_232 : _GEN_4071; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4073 = 3'h6 == pht_windex & 8'he9 == _GEN_14976 ? pht_6_233 : _GEN_4072; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4074 = 3'h6 == pht_windex & 8'hea == _GEN_14976 ? pht_6_234 : _GEN_4073; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4075 = 3'h6 == pht_windex & 8'heb == _GEN_14976 ? pht_6_235 : _GEN_4074; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4076 = 3'h6 == pht_windex & 8'hec == _GEN_14976 ? pht_6_236 : _GEN_4075; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4077 = 3'h6 == pht_windex & 8'hed == _GEN_14976 ? pht_6_237 : _GEN_4076; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4078 = 3'h6 == pht_windex & 8'hee == _GEN_14976 ? pht_6_238 : _GEN_4077; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4079 = 3'h6 == pht_windex & 8'hef == _GEN_14976 ? pht_6_239 : _GEN_4078; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4080 = 3'h6 == pht_windex & 8'hf0 == _GEN_14976 ? pht_6_240 : _GEN_4079; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4081 = 3'h6 == pht_windex & 8'hf1 == _GEN_14976 ? pht_6_241 : _GEN_4080; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4082 = 3'h6 == pht_windex & 8'hf2 == _GEN_14976 ? pht_6_242 : _GEN_4081; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4083 = 3'h6 == pht_windex & 8'hf3 == _GEN_14976 ? pht_6_243 : _GEN_4082; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4084 = 3'h6 == pht_windex & 8'hf4 == _GEN_14976 ? pht_6_244 : _GEN_4083; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4085 = 3'h6 == pht_windex & 8'hf5 == _GEN_14976 ? pht_6_245 : _GEN_4084; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4086 = 3'h6 == pht_windex & 8'hf6 == _GEN_14976 ? pht_6_246 : _GEN_4085; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4087 = 3'h6 == pht_windex & 8'hf7 == _GEN_14976 ? pht_6_247 : _GEN_4086; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4088 = 3'h6 == pht_windex & 8'hf8 == _GEN_14976 ? pht_6_248 : _GEN_4087; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4089 = 3'h6 == pht_windex & 8'hf9 == _GEN_14976 ? pht_6_249 : _GEN_4088; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4090 = 3'h6 == pht_windex & 8'hfa == _GEN_14976 ? pht_6_250 : _GEN_4089; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4091 = 3'h6 == pht_windex & 8'hfb == _GEN_14976 ? pht_6_251 : _GEN_4090; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4092 = 3'h6 == pht_windex & 8'hfc == _GEN_14976 ? pht_6_252 : _GEN_4091; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4093 = 3'h6 == pht_windex & 8'hfd == _GEN_14976 ? pht_6_253 : _GEN_4092; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4094 = 3'h6 == pht_windex & 8'hfe == _GEN_14976 ? pht_6_254 : _GEN_4093; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4095 = 3'h6 == pht_windex & 8'hff == _GEN_14976 ? pht_6_255 : _GEN_4094; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire  _GEN_19584 = 3'h7 == pht_windex; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4096 = 3'h7 == pht_windex & 6'h0 == pht_waddr ? pht_7_0 : _GEN_4095; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4097 = 3'h7 == pht_windex & 6'h1 == pht_waddr ? pht_7_1 : _GEN_4096; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4098 = 3'h7 == pht_windex & 6'h2 == pht_waddr ? pht_7_2 : _GEN_4097; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4099 = 3'h7 == pht_windex & 6'h3 == pht_waddr ? pht_7_3 : _GEN_4098; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4100 = 3'h7 == pht_windex & 6'h4 == pht_waddr ? pht_7_4 : _GEN_4099; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4101 = 3'h7 == pht_windex & 6'h5 == pht_waddr ? pht_7_5 : _GEN_4100; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4102 = 3'h7 == pht_windex & 6'h6 == pht_waddr ? pht_7_6 : _GEN_4101; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4103 = 3'h7 == pht_windex & 6'h7 == pht_waddr ? pht_7_7 : _GEN_4102; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4104 = 3'h7 == pht_windex & 6'h8 == pht_waddr ? pht_7_8 : _GEN_4103; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4105 = 3'h7 == pht_windex & 6'h9 == pht_waddr ? pht_7_9 : _GEN_4104; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4106 = 3'h7 == pht_windex & 6'ha == pht_waddr ? pht_7_10 : _GEN_4105; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4107 = 3'h7 == pht_windex & 6'hb == pht_waddr ? pht_7_11 : _GEN_4106; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4108 = 3'h7 == pht_windex & 6'hc == pht_waddr ? pht_7_12 : _GEN_4107; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4109 = 3'h7 == pht_windex & 6'hd == pht_waddr ? pht_7_13 : _GEN_4108; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4110 = 3'h7 == pht_windex & 6'he == pht_waddr ? pht_7_14 : _GEN_4109; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4111 = 3'h7 == pht_windex & 6'hf == pht_waddr ? pht_7_15 : _GEN_4110; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4112 = 3'h7 == pht_windex & 6'h10 == pht_waddr ? pht_7_16 : _GEN_4111; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4113 = 3'h7 == pht_windex & 6'h11 == pht_waddr ? pht_7_17 : _GEN_4112; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4114 = 3'h7 == pht_windex & 6'h12 == pht_waddr ? pht_7_18 : _GEN_4113; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4115 = 3'h7 == pht_windex & 6'h13 == pht_waddr ? pht_7_19 : _GEN_4114; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4116 = 3'h7 == pht_windex & 6'h14 == pht_waddr ? pht_7_20 : _GEN_4115; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4117 = 3'h7 == pht_windex & 6'h15 == pht_waddr ? pht_7_21 : _GEN_4116; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4118 = 3'h7 == pht_windex & 6'h16 == pht_waddr ? pht_7_22 : _GEN_4117; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4119 = 3'h7 == pht_windex & 6'h17 == pht_waddr ? pht_7_23 : _GEN_4118; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4120 = 3'h7 == pht_windex & 6'h18 == pht_waddr ? pht_7_24 : _GEN_4119; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4121 = 3'h7 == pht_windex & 6'h19 == pht_waddr ? pht_7_25 : _GEN_4120; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4122 = 3'h7 == pht_windex & 6'h1a == pht_waddr ? pht_7_26 : _GEN_4121; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4123 = 3'h7 == pht_windex & 6'h1b == pht_waddr ? pht_7_27 : _GEN_4122; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4124 = 3'h7 == pht_windex & 6'h1c == pht_waddr ? pht_7_28 : _GEN_4123; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4125 = 3'h7 == pht_windex & 6'h1d == pht_waddr ? pht_7_29 : _GEN_4124; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4126 = 3'h7 == pht_windex & 6'h1e == pht_waddr ? pht_7_30 : _GEN_4125; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4127 = 3'h7 == pht_windex & 6'h1f == pht_waddr ? pht_7_31 : _GEN_4126; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4128 = 3'h7 == pht_windex & 6'h20 == pht_waddr ? pht_7_32 : _GEN_4127; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4129 = 3'h7 == pht_windex & 6'h21 == pht_waddr ? pht_7_33 : _GEN_4128; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4130 = 3'h7 == pht_windex & 6'h22 == pht_waddr ? pht_7_34 : _GEN_4129; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4131 = 3'h7 == pht_windex & 6'h23 == pht_waddr ? pht_7_35 : _GEN_4130; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4132 = 3'h7 == pht_windex & 6'h24 == pht_waddr ? pht_7_36 : _GEN_4131; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4133 = 3'h7 == pht_windex & 6'h25 == pht_waddr ? pht_7_37 : _GEN_4132; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4134 = 3'h7 == pht_windex & 6'h26 == pht_waddr ? pht_7_38 : _GEN_4133; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4135 = 3'h7 == pht_windex & 6'h27 == pht_waddr ? pht_7_39 : _GEN_4134; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4136 = 3'h7 == pht_windex & 6'h28 == pht_waddr ? pht_7_40 : _GEN_4135; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4137 = 3'h7 == pht_windex & 6'h29 == pht_waddr ? pht_7_41 : _GEN_4136; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4138 = 3'h7 == pht_windex & 6'h2a == pht_waddr ? pht_7_42 : _GEN_4137; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4139 = 3'h7 == pht_windex & 6'h2b == pht_waddr ? pht_7_43 : _GEN_4138; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4140 = 3'h7 == pht_windex & 6'h2c == pht_waddr ? pht_7_44 : _GEN_4139; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4141 = 3'h7 == pht_windex & 6'h2d == pht_waddr ? pht_7_45 : _GEN_4140; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4142 = 3'h7 == pht_windex & 6'h2e == pht_waddr ? pht_7_46 : _GEN_4141; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4143 = 3'h7 == pht_windex & 6'h2f == pht_waddr ? pht_7_47 : _GEN_4142; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4144 = 3'h7 == pht_windex & 6'h30 == pht_waddr ? pht_7_48 : _GEN_4143; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4145 = 3'h7 == pht_windex & 6'h31 == pht_waddr ? pht_7_49 : _GEN_4144; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4146 = 3'h7 == pht_windex & 6'h32 == pht_waddr ? pht_7_50 : _GEN_4145; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4147 = 3'h7 == pht_windex & 6'h33 == pht_waddr ? pht_7_51 : _GEN_4146; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4148 = 3'h7 == pht_windex & 6'h34 == pht_waddr ? pht_7_52 : _GEN_4147; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4149 = 3'h7 == pht_windex & 6'h35 == pht_waddr ? pht_7_53 : _GEN_4148; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4150 = 3'h7 == pht_windex & 6'h36 == pht_waddr ? pht_7_54 : _GEN_4149; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4151 = 3'h7 == pht_windex & 6'h37 == pht_waddr ? pht_7_55 : _GEN_4150; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4152 = 3'h7 == pht_windex & 6'h38 == pht_waddr ? pht_7_56 : _GEN_4151; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4153 = 3'h7 == pht_windex & 6'h39 == pht_waddr ? pht_7_57 : _GEN_4152; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4154 = 3'h7 == pht_windex & 6'h3a == pht_waddr ? pht_7_58 : _GEN_4153; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4155 = 3'h7 == pht_windex & 6'h3b == pht_waddr ? pht_7_59 : _GEN_4154; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4156 = 3'h7 == pht_windex & 6'h3c == pht_waddr ? pht_7_60 : _GEN_4155; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4157 = 3'h7 == pht_windex & 6'h3d == pht_waddr ? pht_7_61 : _GEN_4156; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4158 = 3'h7 == pht_windex & 6'h3e == pht_waddr ? pht_7_62 : _GEN_4157; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4159 = 3'h7 == pht_windex & 6'h3f == pht_waddr ? pht_7_63 : _GEN_4158; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4160 = 3'h7 == pht_windex & 7'h40 == _GEN_14784 ? pht_7_64 : _GEN_4159; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4161 = 3'h7 == pht_windex & 7'h41 == _GEN_14784 ? pht_7_65 : _GEN_4160; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4162 = 3'h7 == pht_windex & 7'h42 == _GEN_14784 ? pht_7_66 : _GEN_4161; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4163 = 3'h7 == pht_windex & 7'h43 == _GEN_14784 ? pht_7_67 : _GEN_4162; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4164 = 3'h7 == pht_windex & 7'h44 == _GEN_14784 ? pht_7_68 : _GEN_4163; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4165 = 3'h7 == pht_windex & 7'h45 == _GEN_14784 ? pht_7_69 : _GEN_4164; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4166 = 3'h7 == pht_windex & 7'h46 == _GEN_14784 ? pht_7_70 : _GEN_4165; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4167 = 3'h7 == pht_windex & 7'h47 == _GEN_14784 ? pht_7_71 : _GEN_4166; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4168 = 3'h7 == pht_windex & 7'h48 == _GEN_14784 ? pht_7_72 : _GEN_4167; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4169 = 3'h7 == pht_windex & 7'h49 == _GEN_14784 ? pht_7_73 : _GEN_4168; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4170 = 3'h7 == pht_windex & 7'h4a == _GEN_14784 ? pht_7_74 : _GEN_4169; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4171 = 3'h7 == pht_windex & 7'h4b == _GEN_14784 ? pht_7_75 : _GEN_4170; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4172 = 3'h7 == pht_windex & 7'h4c == _GEN_14784 ? pht_7_76 : _GEN_4171; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4173 = 3'h7 == pht_windex & 7'h4d == _GEN_14784 ? pht_7_77 : _GEN_4172; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4174 = 3'h7 == pht_windex & 7'h4e == _GEN_14784 ? pht_7_78 : _GEN_4173; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4175 = 3'h7 == pht_windex & 7'h4f == _GEN_14784 ? pht_7_79 : _GEN_4174; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4176 = 3'h7 == pht_windex & 7'h50 == _GEN_14784 ? pht_7_80 : _GEN_4175; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4177 = 3'h7 == pht_windex & 7'h51 == _GEN_14784 ? pht_7_81 : _GEN_4176; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4178 = 3'h7 == pht_windex & 7'h52 == _GEN_14784 ? pht_7_82 : _GEN_4177; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4179 = 3'h7 == pht_windex & 7'h53 == _GEN_14784 ? pht_7_83 : _GEN_4178; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4180 = 3'h7 == pht_windex & 7'h54 == _GEN_14784 ? pht_7_84 : _GEN_4179; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4181 = 3'h7 == pht_windex & 7'h55 == _GEN_14784 ? pht_7_85 : _GEN_4180; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4182 = 3'h7 == pht_windex & 7'h56 == _GEN_14784 ? pht_7_86 : _GEN_4181; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4183 = 3'h7 == pht_windex & 7'h57 == _GEN_14784 ? pht_7_87 : _GEN_4182; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4184 = 3'h7 == pht_windex & 7'h58 == _GEN_14784 ? pht_7_88 : _GEN_4183; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4185 = 3'h7 == pht_windex & 7'h59 == _GEN_14784 ? pht_7_89 : _GEN_4184; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4186 = 3'h7 == pht_windex & 7'h5a == _GEN_14784 ? pht_7_90 : _GEN_4185; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4187 = 3'h7 == pht_windex & 7'h5b == _GEN_14784 ? pht_7_91 : _GEN_4186; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4188 = 3'h7 == pht_windex & 7'h5c == _GEN_14784 ? pht_7_92 : _GEN_4187; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4189 = 3'h7 == pht_windex & 7'h5d == _GEN_14784 ? pht_7_93 : _GEN_4188; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4190 = 3'h7 == pht_windex & 7'h5e == _GEN_14784 ? pht_7_94 : _GEN_4189; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4191 = 3'h7 == pht_windex & 7'h5f == _GEN_14784 ? pht_7_95 : _GEN_4190; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4192 = 3'h7 == pht_windex & 7'h60 == _GEN_14784 ? pht_7_96 : _GEN_4191; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4193 = 3'h7 == pht_windex & 7'h61 == _GEN_14784 ? pht_7_97 : _GEN_4192; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4194 = 3'h7 == pht_windex & 7'h62 == _GEN_14784 ? pht_7_98 : _GEN_4193; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4195 = 3'h7 == pht_windex & 7'h63 == _GEN_14784 ? pht_7_99 : _GEN_4194; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4196 = 3'h7 == pht_windex & 7'h64 == _GEN_14784 ? pht_7_100 : _GEN_4195; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4197 = 3'h7 == pht_windex & 7'h65 == _GEN_14784 ? pht_7_101 : _GEN_4196; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4198 = 3'h7 == pht_windex & 7'h66 == _GEN_14784 ? pht_7_102 : _GEN_4197; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4199 = 3'h7 == pht_windex & 7'h67 == _GEN_14784 ? pht_7_103 : _GEN_4198; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4200 = 3'h7 == pht_windex & 7'h68 == _GEN_14784 ? pht_7_104 : _GEN_4199; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4201 = 3'h7 == pht_windex & 7'h69 == _GEN_14784 ? pht_7_105 : _GEN_4200; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4202 = 3'h7 == pht_windex & 7'h6a == _GEN_14784 ? pht_7_106 : _GEN_4201; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4203 = 3'h7 == pht_windex & 7'h6b == _GEN_14784 ? pht_7_107 : _GEN_4202; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4204 = 3'h7 == pht_windex & 7'h6c == _GEN_14784 ? pht_7_108 : _GEN_4203; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4205 = 3'h7 == pht_windex & 7'h6d == _GEN_14784 ? pht_7_109 : _GEN_4204; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4206 = 3'h7 == pht_windex & 7'h6e == _GEN_14784 ? pht_7_110 : _GEN_4205; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4207 = 3'h7 == pht_windex & 7'h6f == _GEN_14784 ? pht_7_111 : _GEN_4206; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4208 = 3'h7 == pht_windex & 7'h70 == _GEN_14784 ? pht_7_112 : _GEN_4207; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4209 = 3'h7 == pht_windex & 7'h71 == _GEN_14784 ? pht_7_113 : _GEN_4208; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4210 = 3'h7 == pht_windex & 7'h72 == _GEN_14784 ? pht_7_114 : _GEN_4209; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4211 = 3'h7 == pht_windex & 7'h73 == _GEN_14784 ? pht_7_115 : _GEN_4210; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4212 = 3'h7 == pht_windex & 7'h74 == _GEN_14784 ? pht_7_116 : _GEN_4211; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4213 = 3'h7 == pht_windex & 7'h75 == _GEN_14784 ? pht_7_117 : _GEN_4212; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4214 = 3'h7 == pht_windex & 7'h76 == _GEN_14784 ? pht_7_118 : _GEN_4213; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4215 = 3'h7 == pht_windex & 7'h77 == _GEN_14784 ? pht_7_119 : _GEN_4214; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4216 = 3'h7 == pht_windex & 7'h78 == _GEN_14784 ? pht_7_120 : _GEN_4215; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4217 = 3'h7 == pht_windex & 7'h79 == _GEN_14784 ? pht_7_121 : _GEN_4216; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4218 = 3'h7 == pht_windex & 7'h7a == _GEN_14784 ? pht_7_122 : _GEN_4217; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4219 = 3'h7 == pht_windex & 7'h7b == _GEN_14784 ? pht_7_123 : _GEN_4218; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4220 = 3'h7 == pht_windex & 7'h7c == _GEN_14784 ? pht_7_124 : _GEN_4219; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4221 = 3'h7 == pht_windex & 7'h7d == _GEN_14784 ? pht_7_125 : _GEN_4220; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4222 = 3'h7 == pht_windex & 7'h7e == _GEN_14784 ? pht_7_126 : _GEN_4221; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4223 = 3'h7 == pht_windex & 7'h7f == _GEN_14784 ? pht_7_127 : _GEN_4222; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4224 = 3'h7 == pht_windex & 8'h80 == _GEN_14976 ? pht_7_128 : _GEN_4223; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4225 = 3'h7 == pht_windex & 8'h81 == _GEN_14976 ? pht_7_129 : _GEN_4224; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4226 = 3'h7 == pht_windex & 8'h82 == _GEN_14976 ? pht_7_130 : _GEN_4225; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4227 = 3'h7 == pht_windex & 8'h83 == _GEN_14976 ? pht_7_131 : _GEN_4226; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4228 = 3'h7 == pht_windex & 8'h84 == _GEN_14976 ? pht_7_132 : _GEN_4227; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4229 = 3'h7 == pht_windex & 8'h85 == _GEN_14976 ? pht_7_133 : _GEN_4228; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4230 = 3'h7 == pht_windex & 8'h86 == _GEN_14976 ? pht_7_134 : _GEN_4229; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4231 = 3'h7 == pht_windex & 8'h87 == _GEN_14976 ? pht_7_135 : _GEN_4230; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4232 = 3'h7 == pht_windex & 8'h88 == _GEN_14976 ? pht_7_136 : _GEN_4231; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4233 = 3'h7 == pht_windex & 8'h89 == _GEN_14976 ? pht_7_137 : _GEN_4232; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4234 = 3'h7 == pht_windex & 8'h8a == _GEN_14976 ? pht_7_138 : _GEN_4233; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4235 = 3'h7 == pht_windex & 8'h8b == _GEN_14976 ? pht_7_139 : _GEN_4234; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4236 = 3'h7 == pht_windex & 8'h8c == _GEN_14976 ? pht_7_140 : _GEN_4235; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4237 = 3'h7 == pht_windex & 8'h8d == _GEN_14976 ? pht_7_141 : _GEN_4236; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4238 = 3'h7 == pht_windex & 8'h8e == _GEN_14976 ? pht_7_142 : _GEN_4237; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4239 = 3'h7 == pht_windex & 8'h8f == _GEN_14976 ? pht_7_143 : _GEN_4238; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4240 = 3'h7 == pht_windex & 8'h90 == _GEN_14976 ? pht_7_144 : _GEN_4239; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4241 = 3'h7 == pht_windex & 8'h91 == _GEN_14976 ? pht_7_145 : _GEN_4240; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4242 = 3'h7 == pht_windex & 8'h92 == _GEN_14976 ? pht_7_146 : _GEN_4241; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4243 = 3'h7 == pht_windex & 8'h93 == _GEN_14976 ? pht_7_147 : _GEN_4242; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4244 = 3'h7 == pht_windex & 8'h94 == _GEN_14976 ? pht_7_148 : _GEN_4243; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4245 = 3'h7 == pht_windex & 8'h95 == _GEN_14976 ? pht_7_149 : _GEN_4244; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4246 = 3'h7 == pht_windex & 8'h96 == _GEN_14976 ? pht_7_150 : _GEN_4245; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4247 = 3'h7 == pht_windex & 8'h97 == _GEN_14976 ? pht_7_151 : _GEN_4246; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4248 = 3'h7 == pht_windex & 8'h98 == _GEN_14976 ? pht_7_152 : _GEN_4247; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4249 = 3'h7 == pht_windex & 8'h99 == _GEN_14976 ? pht_7_153 : _GEN_4248; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4250 = 3'h7 == pht_windex & 8'h9a == _GEN_14976 ? pht_7_154 : _GEN_4249; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4251 = 3'h7 == pht_windex & 8'h9b == _GEN_14976 ? pht_7_155 : _GEN_4250; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4252 = 3'h7 == pht_windex & 8'h9c == _GEN_14976 ? pht_7_156 : _GEN_4251; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4253 = 3'h7 == pht_windex & 8'h9d == _GEN_14976 ? pht_7_157 : _GEN_4252; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4254 = 3'h7 == pht_windex & 8'h9e == _GEN_14976 ? pht_7_158 : _GEN_4253; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4255 = 3'h7 == pht_windex & 8'h9f == _GEN_14976 ? pht_7_159 : _GEN_4254; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4256 = 3'h7 == pht_windex & 8'ha0 == _GEN_14976 ? pht_7_160 : _GEN_4255; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4257 = 3'h7 == pht_windex & 8'ha1 == _GEN_14976 ? pht_7_161 : _GEN_4256; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4258 = 3'h7 == pht_windex & 8'ha2 == _GEN_14976 ? pht_7_162 : _GEN_4257; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4259 = 3'h7 == pht_windex & 8'ha3 == _GEN_14976 ? pht_7_163 : _GEN_4258; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4260 = 3'h7 == pht_windex & 8'ha4 == _GEN_14976 ? pht_7_164 : _GEN_4259; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4261 = 3'h7 == pht_windex & 8'ha5 == _GEN_14976 ? pht_7_165 : _GEN_4260; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4262 = 3'h7 == pht_windex & 8'ha6 == _GEN_14976 ? pht_7_166 : _GEN_4261; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4263 = 3'h7 == pht_windex & 8'ha7 == _GEN_14976 ? pht_7_167 : _GEN_4262; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4264 = 3'h7 == pht_windex & 8'ha8 == _GEN_14976 ? pht_7_168 : _GEN_4263; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4265 = 3'h7 == pht_windex & 8'ha9 == _GEN_14976 ? pht_7_169 : _GEN_4264; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4266 = 3'h7 == pht_windex & 8'haa == _GEN_14976 ? pht_7_170 : _GEN_4265; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4267 = 3'h7 == pht_windex & 8'hab == _GEN_14976 ? pht_7_171 : _GEN_4266; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4268 = 3'h7 == pht_windex & 8'hac == _GEN_14976 ? pht_7_172 : _GEN_4267; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4269 = 3'h7 == pht_windex & 8'had == _GEN_14976 ? pht_7_173 : _GEN_4268; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4270 = 3'h7 == pht_windex & 8'hae == _GEN_14976 ? pht_7_174 : _GEN_4269; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4271 = 3'h7 == pht_windex & 8'haf == _GEN_14976 ? pht_7_175 : _GEN_4270; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4272 = 3'h7 == pht_windex & 8'hb0 == _GEN_14976 ? pht_7_176 : _GEN_4271; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4273 = 3'h7 == pht_windex & 8'hb1 == _GEN_14976 ? pht_7_177 : _GEN_4272; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4274 = 3'h7 == pht_windex & 8'hb2 == _GEN_14976 ? pht_7_178 : _GEN_4273; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4275 = 3'h7 == pht_windex & 8'hb3 == _GEN_14976 ? pht_7_179 : _GEN_4274; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4276 = 3'h7 == pht_windex & 8'hb4 == _GEN_14976 ? pht_7_180 : _GEN_4275; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4277 = 3'h7 == pht_windex & 8'hb5 == _GEN_14976 ? pht_7_181 : _GEN_4276; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4278 = 3'h7 == pht_windex & 8'hb6 == _GEN_14976 ? pht_7_182 : _GEN_4277; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4279 = 3'h7 == pht_windex & 8'hb7 == _GEN_14976 ? pht_7_183 : _GEN_4278; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4280 = 3'h7 == pht_windex & 8'hb8 == _GEN_14976 ? pht_7_184 : _GEN_4279; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4281 = 3'h7 == pht_windex & 8'hb9 == _GEN_14976 ? pht_7_185 : _GEN_4280; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4282 = 3'h7 == pht_windex & 8'hba == _GEN_14976 ? pht_7_186 : _GEN_4281; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4283 = 3'h7 == pht_windex & 8'hbb == _GEN_14976 ? pht_7_187 : _GEN_4282; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4284 = 3'h7 == pht_windex & 8'hbc == _GEN_14976 ? pht_7_188 : _GEN_4283; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4285 = 3'h7 == pht_windex & 8'hbd == _GEN_14976 ? pht_7_189 : _GEN_4284; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4286 = 3'h7 == pht_windex & 8'hbe == _GEN_14976 ? pht_7_190 : _GEN_4285; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4287 = 3'h7 == pht_windex & 8'hbf == _GEN_14976 ? pht_7_191 : _GEN_4286; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4288 = 3'h7 == pht_windex & 8'hc0 == _GEN_14976 ? pht_7_192 : _GEN_4287; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4289 = 3'h7 == pht_windex & 8'hc1 == _GEN_14976 ? pht_7_193 : _GEN_4288; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4290 = 3'h7 == pht_windex & 8'hc2 == _GEN_14976 ? pht_7_194 : _GEN_4289; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4291 = 3'h7 == pht_windex & 8'hc3 == _GEN_14976 ? pht_7_195 : _GEN_4290; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4292 = 3'h7 == pht_windex & 8'hc4 == _GEN_14976 ? pht_7_196 : _GEN_4291; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4293 = 3'h7 == pht_windex & 8'hc5 == _GEN_14976 ? pht_7_197 : _GEN_4292; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4294 = 3'h7 == pht_windex & 8'hc6 == _GEN_14976 ? pht_7_198 : _GEN_4293; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4295 = 3'h7 == pht_windex & 8'hc7 == _GEN_14976 ? pht_7_199 : _GEN_4294; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4296 = 3'h7 == pht_windex & 8'hc8 == _GEN_14976 ? pht_7_200 : _GEN_4295; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4297 = 3'h7 == pht_windex & 8'hc9 == _GEN_14976 ? pht_7_201 : _GEN_4296; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4298 = 3'h7 == pht_windex & 8'hca == _GEN_14976 ? pht_7_202 : _GEN_4297; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4299 = 3'h7 == pht_windex & 8'hcb == _GEN_14976 ? pht_7_203 : _GEN_4298; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4300 = 3'h7 == pht_windex & 8'hcc == _GEN_14976 ? pht_7_204 : _GEN_4299; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4301 = 3'h7 == pht_windex & 8'hcd == _GEN_14976 ? pht_7_205 : _GEN_4300; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4302 = 3'h7 == pht_windex & 8'hce == _GEN_14976 ? pht_7_206 : _GEN_4301; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4303 = 3'h7 == pht_windex & 8'hcf == _GEN_14976 ? pht_7_207 : _GEN_4302; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4304 = 3'h7 == pht_windex & 8'hd0 == _GEN_14976 ? pht_7_208 : _GEN_4303; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4305 = 3'h7 == pht_windex & 8'hd1 == _GEN_14976 ? pht_7_209 : _GEN_4304; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4306 = 3'h7 == pht_windex & 8'hd2 == _GEN_14976 ? pht_7_210 : _GEN_4305; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4307 = 3'h7 == pht_windex & 8'hd3 == _GEN_14976 ? pht_7_211 : _GEN_4306; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4308 = 3'h7 == pht_windex & 8'hd4 == _GEN_14976 ? pht_7_212 : _GEN_4307; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4309 = 3'h7 == pht_windex & 8'hd5 == _GEN_14976 ? pht_7_213 : _GEN_4308; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4310 = 3'h7 == pht_windex & 8'hd6 == _GEN_14976 ? pht_7_214 : _GEN_4309; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4311 = 3'h7 == pht_windex & 8'hd7 == _GEN_14976 ? pht_7_215 : _GEN_4310; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4312 = 3'h7 == pht_windex & 8'hd8 == _GEN_14976 ? pht_7_216 : _GEN_4311; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4313 = 3'h7 == pht_windex & 8'hd9 == _GEN_14976 ? pht_7_217 : _GEN_4312; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4314 = 3'h7 == pht_windex & 8'hda == _GEN_14976 ? pht_7_218 : _GEN_4313; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4315 = 3'h7 == pht_windex & 8'hdb == _GEN_14976 ? pht_7_219 : _GEN_4314; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4316 = 3'h7 == pht_windex & 8'hdc == _GEN_14976 ? pht_7_220 : _GEN_4315; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4317 = 3'h7 == pht_windex & 8'hdd == _GEN_14976 ? pht_7_221 : _GEN_4316; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4318 = 3'h7 == pht_windex & 8'hde == _GEN_14976 ? pht_7_222 : _GEN_4317; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4319 = 3'h7 == pht_windex & 8'hdf == _GEN_14976 ? pht_7_223 : _GEN_4318; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4320 = 3'h7 == pht_windex & 8'he0 == _GEN_14976 ? pht_7_224 : _GEN_4319; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4321 = 3'h7 == pht_windex & 8'he1 == _GEN_14976 ? pht_7_225 : _GEN_4320; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4322 = 3'h7 == pht_windex & 8'he2 == _GEN_14976 ? pht_7_226 : _GEN_4321; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4323 = 3'h7 == pht_windex & 8'he3 == _GEN_14976 ? pht_7_227 : _GEN_4322; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4324 = 3'h7 == pht_windex & 8'he4 == _GEN_14976 ? pht_7_228 : _GEN_4323; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4325 = 3'h7 == pht_windex & 8'he5 == _GEN_14976 ? pht_7_229 : _GEN_4324; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4326 = 3'h7 == pht_windex & 8'he6 == _GEN_14976 ? pht_7_230 : _GEN_4325; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4327 = 3'h7 == pht_windex & 8'he7 == _GEN_14976 ? pht_7_231 : _GEN_4326; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4328 = 3'h7 == pht_windex & 8'he8 == _GEN_14976 ? pht_7_232 : _GEN_4327; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4329 = 3'h7 == pht_windex & 8'he9 == _GEN_14976 ? pht_7_233 : _GEN_4328; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4330 = 3'h7 == pht_windex & 8'hea == _GEN_14976 ? pht_7_234 : _GEN_4329; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4331 = 3'h7 == pht_windex & 8'heb == _GEN_14976 ? pht_7_235 : _GEN_4330; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4332 = 3'h7 == pht_windex & 8'hec == _GEN_14976 ? pht_7_236 : _GEN_4331; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4333 = 3'h7 == pht_windex & 8'hed == _GEN_14976 ? pht_7_237 : _GEN_4332; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4334 = 3'h7 == pht_windex & 8'hee == _GEN_14976 ? pht_7_238 : _GEN_4333; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4335 = 3'h7 == pht_windex & 8'hef == _GEN_14976 ? pht_7_239 : _GEN_4334; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4336 = 3'h7 == pht_windex & 8'hf0 == _GEN_14976 ? pht_7_240 : _GEN_4335; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4337 = 3'h7 == pht_windex & 8'hf1 == _GEN_14976 ? pht_7_241 : _GEN_4336; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4338 = 3'h7 == pht_windex & 8'hf2 == _GEN_14976 ? pht_7_242 : _GEN_4337; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4339 = 3'h7 == pht_windex & 8'hf3 == _GEN_14976 ? pht_7_243 : _GEN_4338; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4340 = 3'h7 == pht_windex & 8'hf4 == _GEN_14976 ? pht_7_244 : _GEN_4339; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4341 = 3'h7 == pht_windex & 8'hf5 == _GEN_14976 ? pht_7_245 : _GEN_4340; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4342 = 3'h7 == pht_windex & 8'hf6 == _GEN_14976 ? pht_7_246 : _GEN_4341; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4343 = 3'h7 == pht_windex & 8'hf7 == _GEN_14976 ? pht_7_247 : _GEN_4342; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4344 = 3'h7 == pht_windex & 8'hf8 == _GEN_14976 ? pht_7_248 : _GEN_4343; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4345 = 3'h7 == pht_windex & 8'hf9 == _GEN_14976 ? pht_7_249 : _GEN_4344; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4346 = 3'h7 == pht_windex & 8'hfa == _GEN_14976 ? pht_7_250 : _GEN_4345; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4347 = 3'h7 == pht_windex & 8'hfb == _GEN_14976 ? pht_7_251 : _GEN_4346; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4348 = 3'h7 == pht_windex & 8'hfc == _GEN_14976 ? pht_7_252 : _GEN_4347; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4349 = 3'h7 == pht_windex & 8'hfd == _GEN_14976 ? pht_7_253 : _GEN_4348; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4350 = 3'h7 == pht_windex & 8'hfe == _GEN_14976 ? pht_7_254 : _GEN_4349; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _GEN_4351 = 3'h7 == pht_windex & 8'hff == _GEN_14976 ? pht_7_255 : _GEN_4350; // @[Mux.scala 80:60 Mux.scala 80:60]
  wire [1:0] _pht_T_5 = 2'h1 == _GEN_4351 ? _pht_T_1 : {{1'd0}, io_jmp_packet_jmp}; // @[Mux.scala 80:57]
  wire [1:0] _pht_T_7 = 2'h2 == _GEN_4351 ? _pht_T_2 : _pht_T_5; // @[Mux.scala 80:57]
  reg  btb_0_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_0_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_0_target; // @[BrPredictor.scala 90:20]
  reg  btb_1_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_1_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_1_target; // @[BrPredictor.scala 90:20]
  reg  btb_2_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_2_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_2_target; // @[BrPredictor.scala 90:20]
  reg  btb_3_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_3_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_3_target; // @[BrPredictor.scala 90:20]
  reg  btb_4_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_4_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_4_target; // @[BrPredictor.scala 90:20]
  reg  btb_5_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_5_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_5_target; // @[BrPredictor.scala 90:20]
  reg  btb_6_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_6_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_6_target; // @[BrPredictor.scala 90:20]
  reg  btb_7_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_7_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_7_target; // @[BrPredictor.scala 90:20]
  reg  btb_8_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_8_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_8_target; // @[BrPredictor.scala 90:20]
  reg  btb_9_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_9_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_9_target; // @[BrPredictor.scala 90:20]
  reg  btb_10_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_10_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_10_target; // @[BrPredictor.scala 90:20]
  reg  btb_11_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_11_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_11_target; // @[BrPredictor.scala 90:20]
  reg  btb_12_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_12_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_12_target; // @[BrPredictor.scala 90:20]
  reg  btb_13_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_13_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_13_target; // @[BrPredictor.scala 90:20]
  reg  btb_14_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_14_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_14_target; // @[BrPredictor.scala 90:20]
  reg  btb_15_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_15_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_15_target; // @[BrPredictor.scala 90:20]
  reg  btb_16_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_16_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_16_target; // @[BrPredictor.scala 90:20]
  reg  btb_17_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_17_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_17_target; // @[BrPredictor.scala 90:20]
  reg  btb_18_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_18_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_18_target; // @[BrPredictor.scala 90:20]
  reg  btb_19_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_19_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_19_target; // @[BrPredictor.scala 90:20]
  reg  btb_20_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_20_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_20_target; // @[BrPredictor.scala 90:20]
  reg  btb_21_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_21_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_21_target; // @[BrPredictor.scala 90:20]
  reg  btb_22_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_22_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_22_target; // @[BrPredictor.scala 90:20]
  reg  btb_23_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_23_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_23_target; // @[BrPredictor.scala 90:20]
  reg  btb_24_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_24_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_24_target; // @[BrPredictor.scala 90:20]
  reg  btb_25_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_25_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_25_target; // @[BrPredictor.scala 90:20]
  reg  btb_26_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_26_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_26_target; // @[BrPredictor.scala 90:20]
  reg  btb_27_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_27_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_27_target; // @[BrPredictor.scala 90:20]
  reg  btb_28_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_28_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_28_target; // @[BrPredictor.scala 90:20]
  reg  btb_29_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_29_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_29_target; // @[BrPredictor.scala 90:20]
  reg  btb_30_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_30_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_30_target; // @[BrPredictor.scala 90:20]
  reg  btb_31_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_31_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_31_target; // @[BrPredictor.scala 90:20]
  reg  btb_32_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_32_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_32_target; // @[BrPredictor.scala 90:20]
  reg  btb_33_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_33_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_33_target; // @[BrPredictor.scala 90:20]
  reg  btb_34_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_34_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_34_target; // @[BrPredictor.scala 90:20]
  reg  btb_35_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_35_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_35_target; // @[BrPredictor.scala 90:20]
  reg  btb_36_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_36_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_36_target; // @[BrPredictor.scala 90:20]
  reg  btb_37_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_37_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_37_target; // @[BrPredictor.scala 90:20]
  reg  btb_38_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_38_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_38_target; // @[BrPredictor.scala 90:20]
  reg  btb_39_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_39_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_39_target; // @[BrPredictor.scala 90:20]
  reg  btb_40_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_40_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_40_target; // @[BrPredictor.scala 90:20]
  reg  btb_41_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_41_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_41_target; // @[BrPredictor.scala 90:20]
  reg  btb_42_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_42_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_42_target; // @[BrPredictor.scala 90:20]
  reg  btb_43_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_43_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_43_target; // @[BrPredictor.scala 90:20]
  reg  btb_44_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_44_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_44_target; // @[BrPredictor.scala 90:20]
  reg  btb_45_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_45_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_45_target; // @[BrPredictor.scala 90:20]
  reg  btb_46_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_46_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_46_target; // @[BrPredictor.scala 90:20]
  reg  btb_47_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_47_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_47_target; // @[BrPredictor.scala 90:20]
  reg  btb_48_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_48_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_48_target; // @[BrPredictor.scala 90:20]
  reg  btb_49_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_49_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_49_target; // @[BrPredictor.scala 90:20]
  reg  btb_50_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_50_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_50_target; // @[BrPredictor.scala 90:20]
  reg  btb_51_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_51_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_51_target; // @[BrPredictor.scala 90:20]
  reg  btb_52_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_52_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_52_target; // @[BrPredictor.scala 90:20]
  reg  btb_53_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_53_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_53_target; // @[BrPredictor.scala 90:20]
  reg  btb_54_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_54_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_54_target; // @[BrPredictor.scala 90:20]
  reg  btb_55_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_55_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_55_target; // @[BrPredictor.scala 90:20]
  reg  btb_56_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_56_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_56_target; // @[BrPredictor.scala 90:20]
  reg  btb_57_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_57_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_57_target; // @[BrPredictor.scala 90:20]
  reg  btb_58_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_58_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_58_target; // @[BrPredictor.scala 90:20]
  reg  btb_59_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_59_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_59_target; // @[BrPredictor.scala 90:20]
  reg  btb_60_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_60_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_60_target; // @[BrPredictor.scala 90:20]
  reg  btb_61_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_61_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_61_target; // @[BrPredictor.scala 90:20]
  reg  btb_62_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_62_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_62_target; // @[BrPredictor.scala 90:20]
  reg  btb_63_valid; // @[BrPredictor.scala 90:20]
  reg [7:0] btb_63_tag; // @[BrPredictor.scala 90:20]
  reg [31:0] btb_63_target; // @[BrPredictor.scala 90:20]
  wire [7:0] _GEN_8449 = 6'h1 == bht_raddr ? btb_1_tag : btb_0_tag; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8450 = 6'h2 == bht_raddr ? btb_2_tag : _GEN_8449; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8451 = 6'h3 == bht_raddr ? btb_3_tag : _GEN_8450; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8452 = 6'h4 == bht_raddr ? btb_4_tag : _GEN_8451; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8453 = 6'h5 == bht_raddr ? btb_5_tag : _GEN_8452; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8454 = 6'h6 == bht_raddr ? btb_6_tag : _GEN_8453; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8455 = 6'h7 == bht_raddr ? btb_7_tag : _GEN_8454; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8456 = 6'h8 == bht_raddr ? btb_8_tag : _GEN_8455; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8457 = 6'h9 == bht_raddr ? btb_9_tag : _GEN_8456; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8458 = 6'ha == bht_raddr ? btb_10_tag : _GEN_8457; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8459 = 6'hb == bht_raddr ? btb_11_tag : _GEN_8458; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8460 = 6'hc == bht_raddr ? btb_12_tag : _GEN_8459; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8461 = 6'hd == bht_raddr ? btb_13_tag : _GEN_8460; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8462 = 6'he == bht_raddr ? btb_14_tag : _GEN_8461; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8463 = 6'hf == bht_raddr ? btb_15_tag : _GEN_8462; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8464 = 6'h10 == bht_raddr ? btb_16_tag : _GEN_8463; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8465 = 6'h11 == bht_raddr ? btb_17_tag : _GEN_8464; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8466 = 6'h12 == bht_raddr ? btb_18_tag : _GEN_8465; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8467 = 6'h13 == bht_raddr ? btb_19_tag : _GEN_8466; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8468 = 6'h14 == bht_raddr ? btb_20_tag : _GEN_8467; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8469 = 6'h15 == bht_raddr ? btb_21_tag : _GEN_8468; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8470 = 6'h16 == bht_raddr ? btb_22_tag : _GEN_8469; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8471 = 6'h17 == bht_raddr ? btb_23_tag : _GEN_8470; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8472 = 6'h18 == bht_raddr ? btb_24_tag : _GEN_8471; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8473 = 6'h19 == bht_raddr ? btb_25_tag : _GEN_8472; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8474 = 6'h1a == bht_raddr ? btb_26_tag : _GEN_8473; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8475 = 6'h1b == bht_raddr ? btb_27_tag : _GEN_8474; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8476 = 6'h1c == bht_raddr ? btb_28_tag : _GEN_8475; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8477 = 6'h1d == bht_raddr ? btb_29_tag : _GEN_8476; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8478 = 6'h1e == bht_raddr ? btb_30_tag : _GEN_8477; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8479 = 6'h1f == bht_raddr ? btb_31_tag : _GEN_8478; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8480 = 6'h20 == bht_raddr ? btb_32_tag : _GEN_8479; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8481 = 6'h21 == bht_raddr ? btb_33_tag : _GEN_8480; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8482 = 6'h22 == bht_raddr ? btb_34_tag : _GEN_8481; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8483 = 6'h23 == bht_raddr ? btb_35_tag : _GEN_8482; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8484 = 6'h24 == bht_raddr ? btb_36_tag : _GEN_8483; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8485 = 6'h25 == bht_raddr ? btb_37_tag : _GEN_8484; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8486 = 6'h26 == bht_raddr ? btb_38_tag : _GEN_8485; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8487 = 6'h27 == bht_raddr ? btb_39_tag : _GEN_8486; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8488 = 6'h28 == bht_raddr ? btb_40_tag : _GEN_8487; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8489 = 6'h29 == bht_raddr ? btb_41_tag : _GEN_8488; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8490 = 6'h2a == bht_raddr ? btb_42_tag : _GEN_8489; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8491 = 6'h2b == bht_raddr ? btb_43_tag : _GEN_8490; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8492 = 6'h2c == bht_raddr ? btb_44_tag : _GEN_8491; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8493 = 6'h2d == bht_raddr ? btb_45_tag : _GEN_8492; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8494 = 6'h2e == bht_raddr ? btb_46_tag : _GEN_8493; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8495 = 6'h2f == bht_raddr ? btb_47_tag : _GEN_8494; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8496 = 6'h30 == bht_raddr ? btb_48_tag : _GEN_8495; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8497 = 6'h31 == bht_raddr ? btb_49_tag : _GEN_8496; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8498 = 6'h32 == bht_raddr ? btb_50_tag : _GEN_8497; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8499 = 6'h33 == bht_raddr ? btb_51_tag : _GEN_8498; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8500 = 6'h34 == bht_raddr ? btb_52_tag : _GEN_8499; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8501 = 6'h35 == bht_raddr ? btb_53_tag : _GEN_8500; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8502 = 6'h36 == bht_raddr ? btb_54_tag : _GEN_8501; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8503 = 6'h37 == bht_raddr ? btb_55_tag : _GEN_8502; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8504 = 6'h38 == bht_raddr ? btb_56_tag : _GEN_8503; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8505 = 6'h39 == bht_raddr ? btb_57_tag : _GEN_8504; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8506 = 6'h3a == bht_raddr ? btb_58_tag : _GEN_8505; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8507 = 6'h3b == bht_raddr ? btb_59_tag : _GEN_8506; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8508 = 6'h3c == bht_raddr ? btb_60_tag : _GEN_8507; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8509 = 6'h3d == bht_raddr ? btb_61_tag : _GEN_8508; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8510 = 6'h3e == bht_raddr ? btb_62_tag : _GEN_8509; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire [7:0] _GEN_8511 = 6'h3f == bht_raddr ? btb_63_tag : _GEN_8510; // @[BrPredictor.scala 98:52 BrPredictor.scala 98:52]
  wire  _GEN_8513 = 6'h1 == bht_raddr ? btb_1_valid : btb_0_valid; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8514 = 6'h2 == bht_raddr ? btb_2_valid : _GEN_8513; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8515 = 6'h3 == bht_raddr ? btb_3_valid : _GEN_8514; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8516 = 6'h4 == bht_raddr ? btb_4_valid : _GEN_8515; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8517 = 6'h5 == bht_raddr ? btb_5_valid : _GEN_8516; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8518 = 6'h6 == bht_raddr ? btb_6_valid : _GEN_8517; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8519 = 6'h7 == bht_raddr ? btb_7_valid : _GEN_8518; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8520 = 6'h8 == bht_raddr ? btb_8_valid : _GEN_8519; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8521 = 6'h9 == bht_raddr ? btb_9_valid : _GEN_8520; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8522 = 6'ha == bht_raddr ? btb_10_valid : _GEN_8521; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8523 = 6'hb == bht_raddr ? btb_11_valid : _GEN_8522; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8524 = 6'hc == bht_raddr ? btb_12_valid : _GEN_8523; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8525 = 6'hd == bht_raddr ? btb_13_valid : _GEN_8524; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8526 = 6'he == bht_raddr ? btb_14_valid : _GEN_8525; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8527 = 6'hf == bht_raddr ? btb_15_valid : _GEN_8526; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8528 = 6'h10 == bht_raddr ? btb_16_valid : _GEN_8527; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8529 = 6'h11 == bht_raddr ? btb_17_valid : _GEN_8528; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8530 = 6'h12 == bht_raddr ? btb_18_valid : _GEN_8529; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8531 = 6'h13 == bht_raddr ? btb_19_valid : _GEN_8530; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8532 = 6'h14 == bht_raddr ? btb_20_valid : _GEN_8531; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8533 = 6'h15 == bht_raddr ? btb_21_valid : _GEN_8532; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8534 = 6'h16 == bht_raddr ? btb_22_valid : _GEN_8533; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8535 = 6'h17 == bht_raddr ? btb_23_valid : _GEN_8534; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8536 = 6'h18 == bht_raddr ? btb_24_valid : _GEN_8535; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8537 = 6'h19 == bht_raddr ? btb_25_valid : _GEN_8536; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8538 = 6'h1a == bht_raddr ? btb_26_valid : _GEN_8537; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8539 = 6'h1b == bht_raddr ? btb_27_valid : _GEN_8538; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8540 = 6'h1c == bht_raddr ? btb_28_valid : _GEN_8539; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8541 = 6'h1d == bht_raddr ? btb_29_valid : _GEN_8540; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8542 = 6'h1e == bht_raddr ? btb_30_valid : _GEN_8541; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8543 = 6'h1f == bht_raddr ? btb_31_valid : _GEN_8542; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8544 = 6'h20 == bht_raddr ? btb_32_valid : _GEN_8543; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8545 = 6'h21 == bht_raddr ? btb_33_valid : _GEN_8544; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8546 = 6'h22 == bht_raddr ? btb_34_valid : _GEN_8545; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8547 = 6'h23 == bht_raddr ? btb_35_valid : _GEN_8546; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8548 = 6'h24 == bht_raddr ? btb_36_valid : _GEN_8547; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8549 = 6'h25 == bht_raddr ? btb_37_valid : _GEN_8548; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8550 = 6'h26 == bht_raddr ? btb_38_valid : _GEN_8549; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8551 = 6'h27 == bht_raddr ? btb_39_valid : _GEN_8550; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8552 = 6'h28 == bht_raddr ? btb_40_valid : _GEN_8551; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8553 = 6'h29 == bht_raddr ? btb_41_valid : _GEN_8552; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8554 = 6'h2a == bht_raddr ? btb_42_valid : _GEN_8553; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8555 = 6'h2b == bht_raddr ? btb_43_valid : _GEN_8554; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8556 = 6'h2c == bht_raddr ? btb_44_valid : _GEN_8555; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8557 = 6'h2d == bht_raddr ? btb_45_valid : _GEN_8556; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8558 = 6'h2e == bht_raddr ? btb_46_valid : _GEN_8557; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8559 = 6'h2f == bht_raddr ? btb_47_valid : _GEN_8558; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8560 = 6'h30 == bht_raddr ? btb_48_valid : _GEN_8559; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8561 = 6'h31 == bht_raddr ? btb_49_valid : _GEN_8560; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8562 = 6'h32 == bht_raddr ? btb_50_valid : _GEN_8561; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8563 = 6'h33 == bht_raddr ? btb_51_valid : _GEN_8562; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8564 = 6'h34 == bht_raddr ? btb_52_valid : _GEN_8563; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8565 = 6'h35 == bht_raddr ? btb_53_valid : _GEN_8564; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8566 = 6'h36 == bht_raddr ? btb_54_valid : _GEN_8565; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8567 = 6'h37 == bht_raddr ? btb_55_valid : _GEN_8566; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8568 = 6'h38 == bht_raddr ? btb_56_valid : _GEN_8567; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8569 = 6'h39 == bht_raddr ? btb_57_valid : _GEN_8568; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8570 = 6'h3a == bht_raddr ? btb_58_valid : _GEN_8569; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8571 = 6'h3b == bht_raddr ? btb_59_valid : _GEN_8570; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8572 = 6'h3c == bht_raddr ? btb_60_valid : _GEN_8571; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8573 = 6'h3d == bht_raddr ? btb_61_valid : _GEN_8572; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8574 = 6'h3e == bht_raddr ? btb_62_valid : _GEN_8573; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  _GEN_8575 = 6'h3f == bht_raddr ? btb_63_valid : _GEN_8574; // @[BrPredictor.scala 98:34 BrPredictor.scala 98:34]
  wire  btb_rhit = _GEN_8575 & _GEN_8511 == io_pc[15:8] & io_is_br; // @[BrPredictor.scala 98:68]
  wire  _GEN_8576 = 6'h0 == bht_waddr | btb_0_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8577 = 6'h1 == bht_waddr | btb_1_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8578 = 6'h2 == bht_waddr | btb_2_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8579 = 6'h3 == bht_waddr | btb_3_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8580 = 6'h4 == bht_waddr | btb_4_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8581 = 6'h5 == bht_waddr | btb_5_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8582 = 6'h6 == bht_waddr | btb_6_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8583 = 6'h7 == bht_waddr | btb_7_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8584 = 6'h8 == bht_waddr | btb_8_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8585 = 6'h9 == bht_waddr | btb_9_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8586 = 6'ha == bht_waddr | btb_10_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8587 = 6'hb == bht_waddr | btb_11_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8588 = 6'hc == bht_waddr | btb_12_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8589 = 6'hd == bht_waddr | btb_13_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8590 = 6'he == bht_waddr | btb_14_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8591 = 6'hf == bht_waddr | btb_15_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8592 = 6'h10 == bht_waddr | btb_16_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8593 = 6'h11 == bht_waddr | btb_17_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8594 = 6'h12 == bht_waddr | btb_18_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8595 = 6'h13 == bht_waddr | btb_19_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8596 = 6'h14 == bht_waddr | btb_20_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8597 = 6'h15 == bht_waddr | btb_21_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8598 = 6'h16 == bht_waddr | btb_22_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8599 = 6'h17 == bht_waddr | btb_23_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8600 = 6'h18 == bht_waddr | btb_24_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8601 = 6'h19 == bht_waddr | btb_25_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8602 = 6'h1a == bht_waddr | btb_26_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8603 = 6'h1b == bht_waddr | btb_27_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8604 = 6'h1c == bht_waddr | btb_28_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8605 = 6'h1d == bht_waddr | btb_29_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8606 = 6'h1e == bht_waddr | btb_30_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8607 = 6'h1f == bht_waddr | btb_31_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8608 = 6'h20 == bht_waddr | btb_32_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8609 = 6'h21 == bht_waddr | btb_33_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8610 = 6'h22 == bht_waddr | btb_34_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8611 = 6'h23 == bht_waddr | btb_35_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8612 = 6'h24 == bht_waddr | btb_36_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8613 = 6'h25 == bht_waddr | btb_37_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8614 = 6'h26 == bht_waddr | btb_38_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8615 = 6'h27 == bht_waddr | btb_39_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8616 = 6'h28 == bht_waddr | btb_40_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8617 = 6'h29 == bht_waddr | btb_41_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8618 = 6'h2a == bht_waddr | btb_42_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8619 = 6'h2b == bht_waddr | btb_43_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8620 = 6'h2c == bht_waddr | btb_44_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8621 = 6'h2d == bht_waddr | btb_45_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8622 = 6'h2e == bht_waddr | btb_46_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8623 = 6'h2f == bht_waddr | btb_47_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8624 = 6'h30 == bht_waddr | btb_48_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8625 = 6'h31 == bht_waddr | btb_49_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8626 = 6'h32 == bht_waddr | btb_50_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8627 = 6'h33 == bht_waddr | btb_51_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8628 = 6'h34 == bht_waddr | btb_52_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8629 = 6'h35 == bht_waddr | btb_53_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8630 = 6'h36 == bht_waddr | btb_54_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8631 = 6'h37 == bht_waddr | btb_55_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8632 = 6'h38 == bht_waddr | btb_56_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8633 = 6'h39 == bht_waddr | btb_57_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8634 = 6'h3a == bht_waddr | btb_58_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8635 = 6'h3b == bht_waddr | btb_59_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8636 = 6'h3c == bht_waddr | btb_60_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8637 = 6'h3d == bht_waddr | btb_61_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8638 = 6'h3e == bht_waddr | btb_62_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire  _GEN_8639 = 6'h3f == bht_waddr | btb_63_valid; // @[BrPredictor.scala 104:26 BrPredictor.scala 104:26 BrPredictor.scala 90:20]
  wire [31:0] _pred_pc_T_1 = io_jmp_packet_inst_pc + 32'h4; // @[BrPredictor.scala 111:74]
  wire [31:0] _pred_pc_T_2 = io_jmp_packet_jmp ? io_jmp_packet_jmp_pc : _pred_pc_T_1; // @[BrPredictor.scala 111:19]
  wire [31:0] _GEN_8961 = 6'h1 == bht_raddr ? btb_1_target : btb_0_target; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8962 = 6'h2 == bht_raddr ? btb_2_target : _GEN_8961; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8963 = 6'h3 == bht_raddr ? btb_3_target : _GEN_8962; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8964 = 6'h4 == bht_raddr ? btb_4_target : _GEN_8963; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8965 = 6'h5 == bht_raddr ? btb_5_target : _GEN_8964; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8966 = 6'h6 == bht_raddr ? btb_6_target : _GEN_8965; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8967 = 6'h7 == bht_raddr ? btb_7_target : _GEN_8966; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8968 = 6'h8 == bht_raddr ? btb_8_target : _GEN_8967; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8969 = 6'h9 == bht_raddr ? btb_9_target : _GEN_8968; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8970 = 6'ha == bht_raddr ? btb_10_target : _GEN_8969; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8971 = 6'hb == bht_raddr ? btb_11_target : _GEN_8970; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8972 = 6'hc == bht_raddr ? btb_12_target : _GEN_8971; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8973 = 6'hd == bht_raddr ? btb_13_target : _GEN_8972; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8974 = 6'he == bht_raddr ? btb_14_target : _GEN_8973; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8975 = 6'hf == bht_raddr ? btb_15_target : _GEN_8974; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8976 = 6'h10 == bht_raddr ? btb_16_target : _GEN_8975; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8977 = 6'h11 == bht_raddr ? btb_17_target : _GEN_8976; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8978 = 6'h12 == bht_raddr ? btb_18_target : _GEN_8977; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8979 = 6'h13 == bht_raddr ? btb_19_target : _GEN_8978; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8980 = 6'h14 == bht_raddr ? btb_20_target : _GEN_8979; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8981 = 6'h15 == bht_raddr ? btb_21_target : _GEN_8980; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8982 = 6'h16 == bht_raddr ? btb_22_target : _GEN_8981; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8983 = 6'h17 == bht_raddr ? btb_23_target : _GEN_8982; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8984 = 6'h18 == bht_raddr ? btb_24_target : _GEN_8983; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8985 = 6'h19 == bht_raddr ? btb_25_target : _GEN_8984; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8986 = 6'h1a == bht_raddr ? btb_26_target : _GEN_8985; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8987 = 6'h1b == bht_raddr ? btb_27_target : _GEN_8986; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8988 = 6'h1c == bht_raddr ? btb_28_target : _GEN_8987; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8989 = 6'h1d == bht_raddr ? btb_29_target : _GEN_8988; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8990 = 6'h1e == bht_raddr ? btb_30_target : _GEN_8989; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8991 = 6'h1f == bht_raddr ? btb_31_target : _GEN_8990; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8992 = 6'h20 == bht_raddr ? btb_32_target : _GEN_8991; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8993 = 6'h21 == bht_raddr ? btb_33_target : _GEN_8992; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8994 = 6'h22 == bht_raddr ? btb_34_target : _GEN_8993; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8995 = 6'h23 == bht_raddr ? btb_35_target : _GEN_8994; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8996 = 6'h24 == bht_raddr ? btb_36_target : _GEN_8995; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8997 = 6'h25 == bht_raddr ? btb_37_target : _GEN_8996; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8998 = 6'h26 == bht_raddr ? btb_38_target : _GEN_8997; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_8999 = 6'h27 == bht_raddr ? btb_39_target : _GEN_8998; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9000 = 6'h28 == bht_raddr ? btb_40_target : _GEN_8999; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9001 = 6'h29 == bht_raddr ? btb_41_target : _GEN_9000; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9002 = 6'h2a == bht_raddr ? btb_42_target : _GEN_9001; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9003 = 6'h2b == bht_raddr ? btb_43_target : _GEN_9002; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9004 = 6'h2c == bht_raddr ? btb_44_target : _GEN_9003; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9005 = 6'h2d == bht_raddr ? btb_45_target : _GEN_9004; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9006 = 6'h2e == bht_raddr ? btb_46_target : _GEN_9005; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9007 = 6'h2f == bht_raddr ? btb_47_target : _GEN_9006; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9008 = 6'h30 == bht_raddr ? btb_48_target : _GEN_9007; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9009 = 6'h31 == bht_raddr ? btb_49_target : _GEN_9008; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9010 = 6'h32 == bht_raddr ? btb_50_target : _GEN_9009; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9011 = 6'h33 == bht_raddr ? btb_51_target : _GEN_9010; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9012 = 6'h34 == bht_raddr ? btb_52_target : _GEN_9011; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9013 = 6'h35 == bht_raddr ? btb_53_target : _GEN_9012; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9014 = 6'h36 == bht_raddr ? btb_54_target : _GEN_9013; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9015 = 6'h37 == bht_raddr ? btb_55_target : _GEN_9014; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9016 = 6'h38 == bht_raddr ? btb_56_target : _GEN_9015; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9017 = 6'h39 == bht_raddr ? btb_57_target : _GEN_9016; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9018 = 6'h3a == bht_raddr ? btb_58_target : _GEN_9017; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9019 = 6'h3b == bht_raddr ? btb_59_target : _GEN_9018; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9020 = 6'h3c == bht_raddr ? btb_60_target : _GEN_9019; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9021 = 6'h3d == bht_raddr ? btb_61_target : _GEN_9020; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9022 = 6'h3e == bht_raddr ? btb_62_target : _GEN_9021; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _GEN_9023 = 6'h3f == bht_raddr ? btb_63_target : _GEN_9022; // @[BrPredictor.scala 115:21 BrPredictor.scala 115:21]
  wire [31:0] _pred_pc_T_3 = btb_rhit ? _GEN_9023 : npc; // @[BrPredictor.scala 115:21]
  wire  _GEN_9024 = pht_rdirect & btb_rhit; // @[BrPredictor.scala 113:24 BrPredictor.scala 114:15 BrPredictor.scala 117:15]
  wire [31:0] _GEN_9025 = pht_rdirect ? _pred_pc_T_3 : npc; // @[BrPredictor.scala 113:24 BrPredictor.scala 115:15 BrPredictor.scala 118:15]
  assign io_pred_br = io_jmp_packet_valid & io_jmp_packet_mis ? 1'h0 : _GEN_9024; // @[BrPredictor.scala 109:45 BrPredictor.scala 110:13]
  assign io_pred_pc = io_jmp_packet_valid & io_jmp_packet_mis ? _pred_pc_T_2 : _GEN_9025; // @[BrPredictor.scala 109:45 BrPredictor.scala 111:13]
  always @(posedge clock) begin
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_0 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h0 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_0 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_1 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h1 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_1 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_2 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h2 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_2 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_3 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h3 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_3 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_4 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h4 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_4 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_5 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h5 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_5 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_6 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h6 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_6 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_7 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h7 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_7 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_8 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h8 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_8 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_9 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h9 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_9 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_10 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'ha == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_10 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_11 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'hb == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_11 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_12 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'hc == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_12 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_13 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'hd == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_13 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_14 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'he == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_14 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_15 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'hf == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_15 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_16 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h10 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_16 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_17 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h11 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_17 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_18 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h12 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_18 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_19 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h13 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_19 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_20 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h14 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_20 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_21 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h15 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_21 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_22 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h16 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_22 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_23 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h17 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_23 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_24 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h18 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_24 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_25 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h19 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_25 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_26 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h1a == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_26 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_27 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h1b == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_27 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_28 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h1c == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_28 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_29 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h1d == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_29 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_30 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h1e == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_30 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_31 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h1f == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_31 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_32 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h20 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_32 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_33 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h21 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_33 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_34 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h22 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_34 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_35 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h23 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_35 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_36 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h24 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_36 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_37 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h25 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_37 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_38 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h26 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_38 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_39 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h27 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_39 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_40 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h28 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_40 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_41 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h29 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_41 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_42 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h2a == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_42 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_43 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h2b == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_43 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_44 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h2c == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_44 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_45 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h2d == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_45 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_46 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h2e == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_46 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_47 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h2f == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_47 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_48 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h30 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_48 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_49 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h31 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_49 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_50 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h32 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_50 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_51 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h33 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_51 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_52 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h34 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_52 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_53 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h35 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_53 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_54 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h36 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_54 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_55 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h37 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_55 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_56 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h38 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_56 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_57 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h39 == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_57 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_58 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h3a == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_58 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_59 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h3b == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_59 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_60 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h3c == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_60 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_61 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h3d == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_61 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_62 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h3e == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_62 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 50:20]
      bht_63 <= 6'h0; // @[BrPredictor.scala 50:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 68:27]
      if (6'h3f == bht_waddr) begin // @[BrPredictor.scala 69:20]
        bht_63 <= _bht_T; // @[BrPredictor.scala 69:20]
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_0 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15361) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_0 <= _pht_T_3;
        end else begin
          pht_0_0 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_1 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14659) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_1 <= _pht_T_3;
        end else begin
          pht_0_1 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_2 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14661) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_2 <= _pht_T_3;
        end else begin
          pht_0_2 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_3 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14663) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_3 <= _pht_T_3;
        end else begin
          pht_0_3 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_4 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14665) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_4 <= _pht_T_3;
        end else begin
          pht_0_4 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_5 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14667) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_5 <= _pht_T_3;
        end else begin
          pht_0_5 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_6 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14669) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_6 <= _pht_T_3;
        end else begin
          pht_0_6 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_7 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14671) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_7 <= _pht_T_3;
        end else begin
          pht_0_7 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_8 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14673) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_8 <= _pht_T_3;
        end else begin
          pht_0_8 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_9 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14675) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_9 <= _pht_T_3;
        end else begin
          pht_0_9 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_10 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14677) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_10 <= _pht_T_3;
        end else begin
          pht_0_10 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_11 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14679) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_11 <= _pht_T_3;
        end else begin
          pht_0_11 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_12 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14681) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_12 <= _pht_T_3;
        end else begin
          pht_0_12 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_13 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14683) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_13 <= _pht_T_3;
        end else begin
          pht_0_13 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_14 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14685) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_14 <= _pht_T_3;
        end else begin
          pht_0_14 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_15 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14687) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_15 <= _pht_T_3;
        end else begin
          pht_0_15 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_16 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14689) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_16 <= _pht_T_3;
        end else begin
          pht_0_16 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_17 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14691) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_17 <= _pht_T_3;
        end else begin
          pht_0_17 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_18 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14693) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_18 <= _pht_T_3;
        end else begin
          pht_0_18 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_19 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14695) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_19 <= _pht_T_3;
        end else begin
          pht_0_19 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_20 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14697) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_20 <= _pht_T_3;
        end else begin
          pht_0_20 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_21 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14699) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_21 <= _pht_T_3;
        end else begin
          pht_0_21 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_22 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14701) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_22 <= _pht_T_3;
        end else begin
          pht_0_22 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_23 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14703) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_23 <= _pht_T_3;
        end else begin
          pht_0_23 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_24 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14705) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_24 <= _pht_T_3;
        end else begin
          pht_0_24 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_25 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14707) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_25 <= _pht_T_3;
        end else begin
          pht_0_25 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_26 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14709) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_26 <= _pht_T_3;
        end else begin
          pht_0_26 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_27 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14711) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_27 <= _pht_T_3;
        end else begin
          pht_0_27 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_28 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14713) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_28 <= _pht_T_3;
        end else begin
          pht_0_28 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_29 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14715) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_29 <= _pht_T_3;
        end else begin
          pht_0_29 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_30 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14717) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_30 <= _pht_T_3;
        end else begin
          pht_0_30 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_31 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14719) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_31 <= _pht_T_3;
        end else begin
          pht_0_31 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_32 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14721) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_32 <= _pht_T_3;
        end else begin
          pht_0_32 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_33 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14723) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_33 <= _pht_T_3;
        end else begin
          pht_0_33 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_34 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14725) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_34 <= _pht_T_3;
        end else begin
          pht_0_34 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_35 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14727) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_35 <= _pht_T_3;
        end else begin
          pht_0_35 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_36 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14729) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_36 <= _pht_T_3;
        end else begin
          pht_0_36 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_37 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14731) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_37 <= _pht_T_3;
        end else begin
          pht_0_37 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_38 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14733) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_38 <= _pht_T_3;
        end else begin
          pht_0_38 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_39 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14735) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_39 <= _pht_T_3;
        end else begin
          pht_0_39 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_40 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14737) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_40 <= _pht_T_3;
        end else begin
          pht_0_40 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_41 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14739) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_41 <= _pht_T_3;
        end else begin
          pht_0_41 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_42 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14741) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_42 <= _pht_T_3;
        end else begin
          pht_0_42 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_43 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14743) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_43 <= _pht_T_3;
        end else begin
          pht_0_43 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_44 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14745) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_44 <= _pht_T_3;
        end else begin
          pht_0_44 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_45 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14747) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_45 <= _pht_T_3;
        end else begin
          pht_0_45 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_46 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14749) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_46 <= _pht_T_3;
        end else begin
          pht_0_46 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_47 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14751) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_47 <= _pht_T_3;
        end else begin
          pht_0_47 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_48 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14753) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_48 <= _pht_T_3;
        end else begin
          pht_0_48 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_49 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14755) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_49 <= _pht_T_3;
        end else begin
          pht_0_49 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_50 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14757) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_50 <= _pht_T_3;
        end else begin
          pht_0_50 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_51 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14759) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_51 <= _pht_T_3;
        end else begin
          pht_0_51 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_52 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14761) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_52 <= _pht_T_3;
        end else begin
          pht_0_52 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_53 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14763) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_53 <= _pht_T_3;
        end else begin
          pht_0_53 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_54 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14765) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_54 <= _pht_T_3;
        end else begin
          pht_0_54 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_55 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14767) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_55 <= _pht_T_3;
        end else begin
          pht_0_55 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_56 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14769) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_56 <= _pht_T_3;
        end else begin
          pht_0_56 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_57 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14771) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_57 <= _pht_T_3;
        end else begin
          pht_0_57 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_58 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14773) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_58 <= _pht_T_3;
        end else begin
          pht_0_58 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_59 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14775) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_59 <= _pht_T_3;
        end else begin
          pht_0_59 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_60 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14777) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_60 <= _pht_T_3;
        end else begin
          pht_0_60 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_61 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14779) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_61 <= _pht_T_3;
        end else begin
          pht_0_61 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_62 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14781) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_62 <= _pht_T_3;
        end else begin
          pht_0_62 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_63 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14783) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_63 <= _pht_T_3;
        end else begin
          pht_0_63 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_64 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14786) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_64 <= _pht_T_3;
        end else begin
          pht_0_64 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_65 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14789) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_65 <= _pht_T_3;
        end else begin
          pht_0_65 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_66 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14792) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_66 <= _pht_T_3;
        end else begin
          pht_0_66 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_67 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14795) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_67 <= _pht_T_3;
        end else begin
          pht_0_67 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_68 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14798) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_68 <= _pht_T_3;
        end else begin
          pht_0_68 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_69 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14801) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_69 <= _pht_T_3;
        end else begin
          pht_0_69 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_70 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14804) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_70 <= _pht_T_3;
        end else begin
          pht_0_70 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_71 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14807) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_71 <= _pht_T_3;
        end else begin
          pht_0_71 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_72 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14810) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_72 <= _pht_T_3;
        end else begin
          pht_0_72 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_73 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14813) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_73 <= _pht_T_3;
        end else begin
          pht_0_73 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_74 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14816) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_74 <= _pht_T_3;
        end else begin
          pht_0_74 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_75 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14819) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_75 <= _pht_T_3;
        end else begin
          pht_0_75 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_76 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14822) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_76 <= _pht_T_3;
        end else begin
          pht_0_76 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_77 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14825) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_77 <= _pht_T_3;
        end else begin
          pht_0_77 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_78 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14828) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_78 <= _pht_T_3;
        end else begin
          pht_0_78 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_79 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14831) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_79 <= _pht_T_3;
        end else begin
          pht_0_79 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_80 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14834) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_80 <= _pht_T_3;
        end else begin
          pht_0_80 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_81 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14837) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_81 <= _pht_T_3;
        end else begin
          pht_0_81 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_82 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14840) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_82 <= _pht_T_3;
        end else begin
          pht_0_82 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_83 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14843) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_83 <= _pht_T_3;
        end else begin
          pht_0_83 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_84 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14846) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_84 <= _pht_T_3;
        end else begin
          pht_0_84 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_85 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14849) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_85 <= _pht_T_3;
        end else begin
          pht_0_85 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_86 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14852) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_86 <= _pht_T_3;
        end else begin
          pht_0_86 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_87 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14855) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_87 <= _pht_T_3;
        end else begin
          pht_0_87 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_88 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14858) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_88 <= _pht_T_3;
        end else begin
          pht_0_88 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_89 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14861) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_89 <= _pht_T_3;
        end else begin
          pht_0_89 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_90 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14864) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_90 <= _pht_T_3;
        end else begin
          pht_0_90 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_91 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14867) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_91 <= _pht_T_3;
        end else begin
          pht_0_91 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_92 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14870) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_92 <= _pht_T_3;
        end else begin
          pht_0_92 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_93 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14873) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_93 <= _pht_T_3;
        end else begin
          pht_0_93 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_94 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14876) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_94 <= _pht_T_3;
        end else begin
          pht_0_94 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_95 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14879) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_95 <= _pht_T_3;
        end else begin
          pht_0_95 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_96 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14882) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_96 <= _pht_T_3;
        end else begin
          pht_0_96 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_97 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14885) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_97 <= _pht_T_3;
        end else begin
          pht_0_97 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_98 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14888) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_98 <= _pht_T_3;
        end else begin
          pht_0_98 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_99 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14891) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_99 <= _pht_T_3;
        end else begin
          pht_0_99 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_100 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14894) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_100 <= _pht_T_3;
        end else begin
          pht_0_100 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_101 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14897) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_101 <= _pht_T_3;
        end else begin
          pht_0_101 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_102 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14900) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_102 <= _pht_T_3;
        end else begin
          pht_0_102 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_103 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14903) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_103 <= _pht_T_3;
        end else begin
          pht_0_103 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_104 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14906) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_104 <= _pht_T_3;
        end else begin
          pht_0_104 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_105 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14909) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_105 <= _pht_T_3;
        end else begin
          pht_0_105 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_106 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14912) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_106 <= _pht_T_3;
        end else begin
          pht_0_106 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_107 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14915) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_107 <= _pht_T_3;
        end else begin
          pht_0_107 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_108 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14918) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_108 <= _pht_T_3;
        end else begin
          pht_0_108 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_109 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14921) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_109 <= _pht_T_3;
        end else begin
          pht_0_109 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_110 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14924) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_110 <= _pht_T_3;
        end else begin
          pht_0_110 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_111 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14927) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_111 <= _pht_T_3;
        end else begin
          pht_0_111 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_112 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14930) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_112 <= _pht_T_3;
        end else begin
          pht_0_112 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_113 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14933) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_113 <= _pht_T_3;
        end else begin
          pht_0_113 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_114 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14936) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_114 <= _pht_T_3;
        end else begin
          pht_0_114 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_115 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14939) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_115 <= _pht_T_3;
        end else begin
          pht_0_115 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_116 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14942) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_116 <= _pht_T_3;
        end else begin
          pht_0_116 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_117 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14945) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_117 <= _pht_T_3;
        end else begin
          pht_0_117 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_118 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14948) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_118 <= _pht_T_3;
        end else begin
          pht_0_118 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_119 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14951) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_119 <= _pht_T_3;
        end else begin
          pht_0_119 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_120 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14954) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_120 <= _pht_T_3;
        end else begin
          pht_0_120 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_121 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14957) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_121 <= _pht_T_3;
        end else begin
          pht_0_121 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_122 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14960) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_122 <= _pht_T_3;
        end else begin
          pht_0_122 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_123 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14963) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_123 <= _pht_T_3;
        end else begin
          pht_0_123 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_124 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14966) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_124 <= _pht_T_3;
        end else begin
          pht_0_124 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_125 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14969) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_125 <= _pht_T_3;
        end else begin
          pht_0_125 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_126 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14972) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_126 <= _pht_T_3;
        end else begin
          pht_0_126 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_127 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14975) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_127 <= _pht_T_3;
        end else begin
          pht_0_127 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_128 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14978) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_128 <= _pht_T_3;
        end else begin
          pht_0_128 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_129 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14981) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_129 <= _pht_T_3;
        end else begin
          pht_0_129 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_130 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14984) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_130 <= _pht_T_3;
        end else begin
          pht_0_130 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_131 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14987) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_131 <= _pht_T_3;
        end else begin
          pht_0_131 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_132 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14990) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_132 <= _pht_T_3;
        end else begin
          pht_0_132 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_133 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14993) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_133 <= _pht_T_3;
        end else begin
          pht_0_133 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_134 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14996) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_134 <= _pht_T_3;
        end else begin
          pht_0_134 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_135 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_14999) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_135 <= _pht_T_3;
        end else begin
          pht_0_135 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_136 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15002) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_136 <= _pht_T_3;
        end else begin
          pht_0_136 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_137 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15005) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_137 <= _pht_T_3;
        end else begin
          pht_0_137 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_138 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15008) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_138 <= _pht_T_3;
        end else begin
          pht_0_138 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_139 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15011) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_139 <= _pht_T_3;
        end else begin
          pht_0_139 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_140 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15014) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_140 <= _pht_T_3;
        end else begin
          pht_0_140 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_141 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15017) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_141 <= _pht_T_3;
        end else begin
          pht_0_141 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_142 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15020) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_142 <= _pht_T_3;
        end else begin
          pht_0_142 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_143 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15023) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_143 <= _pht_T_3;
        end else begin
          pht_0_143 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_144 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15026) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_144 <= _pht_T_3;
        end else begin
          pht_0_144 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_145 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15029) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_145 <= _pht_T_3;
        end else begin
          pht_0_145 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_146 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15032) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_146 <= _pht_T_3;
        end else begin
          pht_0_146 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_147 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15035) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_147 <= _pht_T_3;
        end else begin
          pht_0_147 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_148 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15038) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_148 <= _pht_T_3;
        end else begin
          pht_0_148 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_149 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15041) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_149 <= _pht_T_3;
        end else begin
          pht_0_149 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_150 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15044) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_150 <= _pht_T_3;
        end else begin
          pht_0_150 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_151 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15047) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_151 <= _pht_T_3;
        end else begin
          pht_0_151 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_152 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15050) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_152 <= _pht_T_3;
        end else begin
          pht_0_152 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_153 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15053) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_153 <= _pht_T_3;
        end else begin
          pht_0_153 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_154 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15056) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_154 <= _pht_T_3;
        end else begin
          pht_0_154 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_155 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15059) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_155 <= _pht_T_3;
        end else begin
          pht_0_155 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_156 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15062) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_156 <= _pht_T_3;
        end else begin
          pht_0_156 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_157 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15065) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_157 <= _pht_T_3;
        end else begin
          pht_0_157 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_158 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15068) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_158 <= _pht_T_3;
        end else begin
          pht_0_158 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_159 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15071) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_159 <= _pht_T_3;
        end else begin
          pht_0_159 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_160 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15074) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_160 <= _pht_T_3;
        end else begin
          pht_0_160 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_161 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15077) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_161 <= _pht_T_3;
        end else begin
          pht_0_161 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_162 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15080) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_162 <= _pht_T_3;
        end else begin
          pht_0_162 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_163 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15083) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_163 <= _pht_T_3;
        end else begin
          pht_0_163 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_164 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15086) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_164 <= _pht_T_3;
        end else begin
          pht_0_164 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_165 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15089) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_165 <= _pht_T_3;
        end else begin
          pht_0_165 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_166 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15092) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_166 <= _pht_T_3;
        end else begin
          pht_0_166 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_167 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15095) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_167 <= _pht_T_3;
        end else begin
          pht_0_167 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_168 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15098) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_168 <= _pht_T_3;
        end else begin
          pht_0_168 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_169 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15101) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_169 <= _pht_T_3;
        end else begin
          pht_0_169 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_170 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15104) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_170 <= _pht_T_3;
        end else begin
          pht_0_170 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_171 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15107) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_171 <= _pht_T_3;
        end else begin
          pht_0_171 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_172 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15110) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_172 <= _pht_T_3;
        end else begin
          pht_0_172 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_173 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15113) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_173 <= _pht_T_3;
        end else begin
          pht_0_173 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_174 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15116) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_174 <= _pht_T_3;
        end else begin
          pht_0_174 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_175 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15119) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_175 <= _pht_T_3;
        end else begin
          pht_0_175 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_176 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15122) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_176 <= _pht_T_3;
        end else begin
          pht_0_176 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_177 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15125) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_177 <= _pht_T_3;
        end else begin
          pht_0_177 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_178 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15128) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_178 <= _pht_T_3;
        end else begin
          pht_0_178 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_179 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15131) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_179 <= _pht_T_3;
        end else begin
          pht_0_179 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_180 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15134) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_180 <= _pht_T_3;
        end else begin
          pht_0_180 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_181 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15137) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_181 <= _pht_T_3;
        end else begin
          pht_0_181 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_182 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15140) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_182 <= _pht_T_3;
        end else begin
          pht_0_182 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_183 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15143) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_183 <= _pht_T_3;
        end else begin
          pht_0_183 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_184 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15146) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_184 <= _pht_T_3;
        end else begin
          pht_0_184 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_185 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15149) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_185 <= _pht_T_3;
        end else begin
          pht_0_185 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_186 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15152) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_186 <= _pht_T_3;
        end else begin
          pht_0_186 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_187 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15155) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_187 <= _pht_T_3;
        end else begin
          pht_0_187 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_188 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15158) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_188 <= _pht_T_3;
        end else begin
          pht_0_188 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_189 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15161) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_189 <= _pht_T_3;
        end else begin
          pht_0_189 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_190 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15164) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_190 <= _pht_T_3;
        end else begin
          pht_0_190 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_191 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15167) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_191 <= _pht_T_3;
        end else begin
          pht_0_191 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_192 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15170) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_192 <= _pht_T_3;
        end else begin
          pht_0_192 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_193 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15173) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_193 <= _pht_T_3;
        end else begin
          pht_0_193 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_194 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15176) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_194 <= _pht_T_3;
        end else begin
          pht_0_194 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_195 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15179) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_195 <= _pht_T_3;
        end else begin
          pht_0_195 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_196 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15182) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_196 <= _pht_T_3;
        end else begin
          pht_0_196 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_197 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15185) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_197 <= _pht_T_3;
        end else begin
          pht_0_197 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_198 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15188) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_198 <= _pht_T_3;
        end else begin
          pht_0_198 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_199 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15191) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_199 <= _pht_T_3;
        end else begin
          pht_0_199 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_200 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15194) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_200 <= _pht_T_3;
        end else begin
          pht_0_200 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_201 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15197) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_201 <= _pht_T_3;
        end else begin
          pht_0_201 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_202 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15200) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_202 <= _pht_T_3;
        end else begin
          pht_0_202 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_203 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15203) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_203 <= _pht_T_3;
        end else begin
          pht_0_203 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_204 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15206) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_204 <= _pht_T_3;
        end else begin
          pht_0_204 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_205 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15209) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_205 <= _pht_T_3;
        end else begin
          pht_0_205 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_206 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15212) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_206 <= _pht_T_3;
        end else begin
          pht_0_206 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_207 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15215) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_207 <= _pht_T_3;
        end else begin
          pht_0_207 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_208 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15218) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_208 <= _pht_T_3;
        end else begin
          pht_0_208 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_209 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15221) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_209 <= _pht_T_3;
        end else begin
          pht_0_209 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_210 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15224) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_210 <= _pht_T_3;
        end else begin
          pht_0_210 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_211 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15227) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_211 <= _pht_T_3;
        end else begin
          pht_0_211 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_212 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15230) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_212 <= _pht_T_3;
        end else begin
          pht_0_212 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_213 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15233) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_213 <= _pht_T_3;
        end else begin
          pht_0_213 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_214 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15236) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_214 <= _pht_T_3;
        end else begin
          pht_0_214 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_215 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15239) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_215 <= _pht_T_3;
        end else begin
          pht_0_215 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_216 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15242) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_216 <= _pht_T_3;
        end else begin
          pht_0_216 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_217 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15245) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_217 <= _pht_T_3;
        end else begin
          pht_0_217 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_218 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15248) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_218 <= _pht_T_3;
        end else begin
          pht_0_218 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_219 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15251) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_219 <= _pht_T_3;
        end else begin
          pht_0_219 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_220 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15254) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_220 <= _pht_T_3;
        end else begin
          pht_0_220 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_221 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15257) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_221 <= _pht_T_3;
        end else begin
          pht_0_221 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_222 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15260) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_222 <= _pht_T_3;
        end else begin
          pht_0_222 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_223 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15263) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_223 <= _pht_T_3;
        end else begin
          pht_0_223 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_224 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15266) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_224 <= _pht_T_3;
        end else begin
          pht_0_224 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_225 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15269) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_225 <= _pht_T_3;
        end else begin
          pht_0_225 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_226 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15272) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_226 <= _pht_T_3;
        end else begin
          pht_0_226 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_227 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15275) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_227 <= _pht_T_3;
        end else begin
          pht_0_227 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_228 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15278) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_228 <= _pht_T_3;
        end else begin
          pht_0_228 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_229 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15281) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_229 <= _pht_T_3;
        end else begin
          pht_0_229 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_230 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15284) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_230 <= _pht_T_3;
        end else begin
          pht_0_230 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_231 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15287) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_231 <= _pht_T_3;
        end else begin
          pht_0_231 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_232 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15290) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_232 <= _pht_T_3;
        end else begin
          pht_0_232 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_233 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15293) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_233 <= _pht_T_3;
        end else begin
          pht_0_233 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_234 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15296) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_234 <= _pht_T_3;
        end else begin
          pht_0_234 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_235 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15299) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_235 <= _pht_T_3;
        end else begin
          pht_0_235 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_236 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15302) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_236 <= _pht_T_3;
        end else begin
          pht_0_236 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_237 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15305) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_237 <= _pht_T_3;
        end else begin
          pht_0_237 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_238 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15308) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_238 <= _pht_T_3;
        end else begin
          pht_0_238 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_239 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15311) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_239 <= _pht_T_3;
        end else begin
          pht_0_239 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_240 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15314) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_240 <= _pht_T_3;
        end else begin
          pht_0_240 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_241 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15317) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_241 <= _pht_T_3;
        end else begin
          pht_0_241 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_242 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15320) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_242 <= _pht_T_3;
        end else begin
          pht_0_242 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_243 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15323) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_243 <= _pht_T_3;
        end else begin
          pht_0_243 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_244 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15326) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_244 <= _pht_T_3;
        end else begin
          pht_0_244 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_245 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15329) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_245 <= _pht_T_3;
        end else begin
          pht_0_245 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_246 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15332) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_246 <= _pht_T_3;
        end else begin
          pht_0_246 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_247 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15335) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_247 <= _pht_T_3;
        end else begin
          pht_0_247 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_248 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15338) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_248 <= _pht_T_3;
        end else begin
          pht_0_248 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_249 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15341) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_249 <= _pht_T_3;
        end else begin
          pht_0_249 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_250 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15344) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_250 <= _pht_T_3;
        end else begin
          pht_0_250 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_251 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15347) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_251 <= _pht_T_3;
        end else begin
          pht_0_251 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_252 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15350) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_252 <= _pht_T_3;
        end else begin
          pht_0_252 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_253 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15353) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_253 <= _pht_T_3;
        end else begin
          pht_0_253 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_254 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15356) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_254 <= _pht_T_3;
        end else begin
          pht_0_254 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_0_255 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_14658 & _GEN_15359) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_0_255 <= _pht_T_3;
        end else begin
          pht_0_255 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_0 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15361) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_0 <= _pht_T_3;
        end else begin
          pht_1_0 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_1 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14659) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_1 <= _pht_T_3;
        end else begin
          pht_1_1 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_2 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14661) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_2 <= _pht_T_3;
        end else begin
          pht_1_2 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_3 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14663) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_3 <= _pht_T_3;
        end else begin
          pht_1_3 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_4 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14665) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_4 <= _pht_T_3;
        end else begin
          pht_1_4 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_5 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14667) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_5 <= _pht_T_3;
        end else begin
          pht_1_5 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_6 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14669) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_6 <= _pht_T_3;
        end else begin
          pht_1_6 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_7 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14671) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_7 <= _pht_T_3;
        end else begin
          pht_1_7 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_8 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14673) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_8 <= _pht_T_3;
        end else begin
          pht_1_8 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_9 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14675) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_9 <= _pht_T_3;
        end else begin
          pht_1_9 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_10 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14677) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_10 <= _pht_T_3;
        end else begin
          pht_1_10 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_11 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14679) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_11 <= _pht_T_3;
        end else begin
          pht_1_11 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_12 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14681) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_12 <= _pht_T_3;
        end else begin
          pht_1_12 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_13 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14683) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_13 <= _pht_T_3;
        end else begin
          pht_1_13 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_14 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14685) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_14 <= _pht_T_3;
        end else begin
          pht_1_14 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_15 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14687) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_15 <= _pht_T_3;
        end else begin
          pht_1_15 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_16 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14689) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_16 <= _pht_T_3;
        end else begin
          pht_1_16 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_17 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14691) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_17 <= _pht_T_3;
        end else begin
          pht_1_17 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_18 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14693) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_18 <= _pht_T_3;
        end else begin
          pht_1_18 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_19 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14695) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_19 <= _pht_T_3;
        end else begin
          pht_1_19 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_20 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14697) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_20 <= _pht_T_3;
        end else begin
          pht_1_20 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_21 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14699) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_21 <= _pht_T_3;
        end else begin
          pht_1_21 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_22 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14701) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_22 <= _pht_T_3;
        end else begin
          pht_1_22 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_23 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14703) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_23 <= _pht_T_3;
        end else begin
          pht_1_23 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_24 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14705) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_24 <= _pht_T_3;
        end else begin
          pht_1_24 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_25 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14707) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_25 <= _pht_T_3;
        end else begin
          pht_1_25 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_26 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14709) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_26 <= _pht_T_3;
        end else begin
          pht_1_26 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_27 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14711) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_27 <= _pht_T_3;
        end else begin
          pht_1_27 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_28 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14713) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_28 <= _pht_T_3;
        end else begin
          pht_1_28 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_29 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14715) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_29 <= _pht_T_3;
        end else begin
          pht_1_29 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_30 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14717) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_30 <= _pht_T_3;
        end else begin
          pht_1_30 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_31 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14719) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_31 <= _pht_T_3;
        end else begin
          pht_1_31 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_32 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14721) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_32 <= _pht_T_3;
        end else begin
          pht_1_32 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_33 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14723) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_33 <= _pht_T_3;
        end else begin
          pht_1_33 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_34 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14725) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_34 <= _pht_T_3;
        end else begin
          pht_1_34 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_35 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14727) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_35 <= _pht_T_3;
        end else begin
          pht_1_35 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_36 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14729) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_36 <= _pht_T_3;
        end else begin
          pht_1_36 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_37 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14731) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_37 <= _pht_T_3;
        end else begin
          pht_1_37 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_38 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14733) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_38 <= _pht_T_3;
        end else begin
          pht_1_38 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_39 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14735) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_39 <= _pht_T_3;
        end else begin
          pht_1_39 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_40 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14737) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_40 <= _pht_T_3;
        end else begin
          pht_1_40 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_41 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14739) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_41 <= _pht_T_3;
        end else begin
          pht_1_41 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_42 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14741) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_42 <= _pht_T_3;
        end else begin
          pht_1_42 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_43 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14743) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_43 <= _pht_T_3;
        end else begin
          pht_1_43 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_44 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14745) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_44 <= _pht_T_3;
        end else begin
          pht_1_44 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_45 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14747) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_45 <= _pht_T_3;
        end else begin
          pht_1_45 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_46 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14749) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_46 <= _pht_T_3;
        end else begin
          pht_1_46 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_47 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14751) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_47 <= _pht_T_3;
        end else begin
          pht_1_47 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_48 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14753) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_48 <= _pht_T_3;
        end else begin
          pht_1_48 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_49 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14755) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_49 <= _pht_T_3;
        end else begin
          pht_1_49 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_50 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14757) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_50 <= _pht_T_3;
        end else begin
          pht_1_50 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_51 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14759) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_51 <= _pht_T_3;
        end else begin
          pht_1_51 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_52 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14761) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_52 <= _pht_T_3;
        end else begin
          pht_1_52 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_53 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14763) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_53 <= _pht_T_3;
        end else begin
          pht_1_53 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_54 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14765) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_54 <= _pht_T_3;
        end else begin
          pht_1_54 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_55 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14767) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_55 <= _pht_T_3;
        end else begin
          pht_1_55 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_56 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14769) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_56 <= _pht_T_3;
        end else begin
          pht_1_56 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_57 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14771) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_57 <= _pht_T_3;
        end else begin
          pht_1_57 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_58 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14773) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_58 <= _pht_T_3;
        end else begin
          pht_1_58 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_59 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14775) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_59 <= _pht_T_3;
        end else begin
          pht_1_59 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_60 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14777) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_60 <= _pht_T_3;
        end else begin
          pht_1_60 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_61 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14779) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_61 <= _pht_T_3;
        end else begin
          pht_1_61 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_62 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14781) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_62 <= _pht_T_3;
        end else begin
          pht_1_62 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_63 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14783) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_63 <= _pht_T_3;
        end else begin
          pht_1_63 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_64 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14786) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_64 <= _pht_T_3;
        end else begin
          pht_1_64 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_65 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14789) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_65 <= _pht_T_3;
        end else begin
          pht_1_65 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_66 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14792) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_66 <= _pht_T_3;
        end else begin
          pht_1_66 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_67 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14795) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_67 <= _pht_T_3;
        end else begin
          pht_1_67 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_68 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14798) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_68 <= _pht_T_3;
        end else begin
          pht_1_68 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_69 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14801) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_69 <= _pht_T_3;
        end else begin
          pht_1_69 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_70 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14804) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_70 <= _pht_T_3;
        end else begin
          pht_1_70 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_71 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14807) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_71 <= _pht_T_3;
        end else begin
          pht_1_71 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_72 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14810) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_72 <= _pht_T_3;
        end else begin
          pht_1_72 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_73 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14813) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_73 <= _pht_T_3;
        end else begin
          pht_1_73 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_74 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14816) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_74 <= _pht_T_3;
        end else begin
          pht_1_74 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_75 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14819) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_75 <= _pht_T_3;
        end else begin
          pht_1_75 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_76 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14822) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_76 <= _pht_T_3;
        end else begin
          pht_1_76 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_77 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14825) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_77 <= _pht_T_3;
        end else begin
          pht_1_77 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_78 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14828) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_78 <= _pht_T_3;
        end else begin
          pht_1_78 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_79 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14831) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_79 <= _pht_T_3;
        end else begin
          pht_1_79 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_80 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14834) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_80 <= _pht_T_3;
        end else begin
          pht_1_80 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_81 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14837) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_81 <= _pht_T_3;
        end else begin
          pht_1_81 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_82 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14840) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_82 <= _pht_T_3;
        end else begin
          pht_1_82 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_83 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14843) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_83 <= _pht_T_3;
        end else begin
          pht_1_83 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_84 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14846) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_84 <= _pht_T_3;
        end else begin
          pht_1_84 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_85 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14849) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_85 <= _pht_T_3;
        end else begin
          pht_1_85 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_86 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14852) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_86 <= _pht_T_3;
        end else begin
          pht_1_86 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_87 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14855) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_87 <= _pht_T_3;
        end else begin
          pht_1_87 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_88 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14858) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_88 <= _pht_T_3;
        end else begin
          pht_1_88 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_89 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14861) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_89 <= _pht_T_3;
        end else begin
          pht_1_89 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_90 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14864) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_90 <= _pht_T_3;
        end else begin
          pht_1_90 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_91 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14867) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_91 <= _pht_T_3;
        end else begin
          pht_1_91 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_92 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14870) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_92 <= _pht_T_3;
        end else begin
          pht_1_92 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_93 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14873) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_93 <= _pht_T_3;
        end else begin
          pht_1_93 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_94 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14876) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_94 <= _pht_T_3;
        end else begin
          pht_1_94 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_95 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14879) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_95 <= _pht_T_3;
        end else begin
          pht_1_95 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_96 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14882) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_96 <= _pht_T_3;
        end else begin
          pht_1_96 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_97 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14885) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_97 <= _pht_T_3;
        end else begin
          pht_1_97 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_98 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14888) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_98 <= _pht_T_3;
        end else begin
          pht_1_98 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_99 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14891) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_99 <= _pht_T_3;
        end else begin
          pht_1_99 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_100 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14894) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_100 <= _pht_T_3;
        end else begin
          pht_1_100 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_101 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14897) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_101 <= _pht_T_3;
        end else begin
          pht_1_101 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_102 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14900) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_102 <= _pht_T_3;
        end else begin
          pht_1_102 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_103 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14903) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_103 <= _pht_T_3;
        end else begin
          pht_1_103 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_104 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14906) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_104 <= _pht_T_3;
        end else begin
          pht_1_104 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_105 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14909) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_105 <= _pht_T_3;
        end else begin
          pht_1_105 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_106 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14912) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_106 <= _pht_T_3;
        end else begin
          pht_1_106 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_107 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14915) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_107 <= _pht_T_3;
        end else begin
          pht_1_107 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_108 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14918) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_108 <= _pht_T_3;
        end else begin
          pht_1_108 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_109 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14921) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_109 <= _pht_T_3;
        end else begin
          pht_1_109 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_110 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14924) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_110 <= _pht_T_3;
        end else begin
          pht_1_110 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_111 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14927) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_111 <= _pht_T_3;
        end else begin
          pht_1_111 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_112 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14930) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_112 <= _pht_T_3;
        end else begin
          pht_1_112 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_113 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14933) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_113 <= _pht_T_3;
        end else begin
          pht_1_113 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_114 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14936) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_114 <= _pht_T_3;
        end else begin
          pht_1_114 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_115 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14939) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_115 <= _pht_T_3;
        end else begin
          pht_1_115 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_116 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14942) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_116 <= _pht_T_3;
        end else begin
          pht_1_116 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_117 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14945) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_117 <= _pht_T_3;
        end else begin
          pht_1_117 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_118 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14948) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_118 <= _pht_T_3;
        end else begin
          pht_1_118 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_119 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14951) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_119 <= _pht_T_3;
        end else begin
          pht_1_119 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_120 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14954) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_120 <= _pht_T_3;
        end else begin
          pht_1_120 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_121 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14957) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_121 <= _pht_T_3;
        end else begin
          pht_1_121 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_122 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14960) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_122 <= _pht_T_3;
        end else begin
          pht_1_122 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_123 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14963) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_123 <= _pht_T_3;
        end else begin
          pht_1_123 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_124 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14966) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_124 <= _pht_T_3;
        end else begin
          pht_1_124 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_125 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14969) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_125 <= _pht_T_3;
        end else begin
          pht_1_125 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_126 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14972) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_126 <= _pht_T_3;
        end else begin
          pht_1_126 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_127 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14975) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_127 <= _pht_T_3;
        end else begin
          pht_1_127 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_128 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14978) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_128 <= _pht_T_3;
        end else begin
          pht_1_128 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_129 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14981) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_129 <= _pht_T_3;
        end else begin
          pht_1_129 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_130 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14984) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_130 <= _pht_T_3;
        end else begin
          pht_1_130 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_131 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14987) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_131 <= _pht_T_3;
        end else begin
          pht_1_131 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_132 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14990) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_132 <= _pht_T_3;
        end else begin
          pht_1_132 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_133 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14993) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_133 <= _pht_T_3;
        end else begin
          pht_1_133 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_134 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14996) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_134 <= _pht_T_3;
        end else begin
          pht_1_134 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_135 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_14999) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_135 <= _pht_T_3;
        end else begin
          pht_1_135 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_136 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15002) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_136 <= _pht_T_3;
        end else begin
          pht_1_136 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_137 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15005) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_137 <= _pht_T_3;
        end else begin
          pht_1_137 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_138 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15008) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_138 <= _pht_T_3;
        end else begin
          pht_1_138 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_139 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15011) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_139 <= _pht_T_3;
        end else begin
          pht_1_139 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_140 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15014) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_140 <= _pht_T_3;
        end else begin
          pht_1_140 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_141 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15017) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_141 <= _pht_T_3;
        end else begin
          pht_1_141 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_142 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15020) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_142 <= _pht_T_3;
        end else begin
          pht_1_142 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_143 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15023) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_143 <= _pht_T_3;
        end else begin
          pht_1_143 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_144 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15026) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_144 <= _pht_T_3;
        end else begin
          pht_1_144 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_145 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15029) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_145 <= _pht_T_3;
        end else begin
          pht_1_145 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_146 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15032) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_146 <= _pht_T_3;
        end else begin
          pht_1_146 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_147 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15035) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_147 <= _pht_T_3;
        end else begin
          pht_1_147 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_148 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15038) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_148 <= _pht_T_3;
        end else begin
          pht_1_148 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_149 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15041) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_149 <= _pht_T_3;
        end else begin
          pht_1_149 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_150 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15044) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_150 <= _pht_T_3;
        end else begin
          pht_1_150 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_151 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15047) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_151 <= _pht_T_3;
        end else begin
          pht_1_151 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_152 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15050) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_152 <= _pht_T_3;
        end else begin
          pht_1_152 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_153 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15053) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_153 <= _pht_T_3;
        end else begin
          pht_1_153 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_154 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15056) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_154 <= _pht_T_3;
        end else begin
          pht_1_154 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_155 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15059) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_155 <= _pht_T_3;
        end else begin
          pht_1_155 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_156 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15062) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_156 <= _pht_T_3;
        end else begin
          pht_1_156 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_157 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15065) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_157 <= _pht_T_3;
        end else begin
          pht_1_157 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_158 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15068) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_158 <= _pht_T_3;
        end else begin
          pht_1_158 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_159 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15071) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_159 <= _pht_T_3;
        end else begin
          pht_1_159 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_160 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15074) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_160 <= _pht_T_3;
        end else begin
          pht_1_160 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_161 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15077) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_161 <= _pht_T_3;
        end else begin
          pht_1_161 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_162 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15080) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_162 <= _pht_T_3;
        end else begin
          pht_1_162 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_163 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15083) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_163 <= _pht_T_3;
        end else begin
          pht_1_163 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_164 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15086) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_164 <= _pht_T_3;
        end else begin
          pht_1_164 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_165 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15089) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_165 <= _pht_T_3;
        end else begin
          pht_1_165 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_166 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15092) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_166 <= _pht_T_3;
        end else begin
          pht_1_166 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_167 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15095) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_167 <= _pht_T_3;
        end else begin
          pht_1_167 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_168 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15098) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_168 <= _pht_T_3;
        end else begin
          pht_1_168 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_169 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15101) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_169 <= _pht_T_3;
        end else begin
          pht_1_169 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_170 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15104) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_170 <= _pht_T_3;
        end else begin
          pht_1_170 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_171 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15107) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_171 <= _pht_T_3;
        end else begin
          pht_1_171 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_172 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15110) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_172 <= _pht_T_3;
        end else begin
          pht_1_172 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_173 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15113) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_173 <= _pht_T_3;
        end else begin
          pht_1_173 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_174 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15116) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_174 <= _pht_T_3;
        end else begin
          pht_1_174 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_175 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15119) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_175 <= _pht_T_3;
        end else begin
          pht_1_175 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_176 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15122) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_176 <= _pht_T_3;
        end else begin
          pht_1_176 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_177 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15125) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_177 <= _pht_T_3;
        end else begin
          pht_1_177 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_178 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15128) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_178 <= _pht_T_3;
        end else begin
          pht_1_178 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_179 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15131) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_179 <= _pht_T_3;
        end else begin
          pht_1_179 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_180 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15134) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_180 <= _pht_T_3;
        end else begin
          pht_1_180 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_181 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15137) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_181 <= _pht_T_3;
        end else begin
          pht_1_181 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_182 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15140) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_182 <= _pht_T_3;
        end else begin
          pht_1_182 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_183 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15143) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_183 <= _pht_T_3;
        end else begin
          pht_1_183 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_184 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15146) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_184 <= _pht_T_3;
        end else begin
          pht_1_184 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_185 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15149) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_185 <= _pht_T_3;
        end else begin
          pht_1_185 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_186 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15152) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_186 <= _pht_T_3;
        end else begin
          pht_1_186 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_187 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15155) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_187 <= _pht_T_3;
        end else begin
          pht_1_187 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_188 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15158) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_188 <= _pht_T_3;
        end else begin
          pht_1_188 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_189 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15161) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_189 <= _pht_T_3;
        end else begin
          pht_1_189 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_190 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15164) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_190 <= _pht_T_3;
        end else begin
          pht_1_190 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_191 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15167) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_191 <= _pht_T_3;
        end else begin
          pht_1_191 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_192 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15170) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_192 <= _pht_T_3;
        end else begin
          pht_1_192 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_193 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15173) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_193 <= _pht_T_3;
        end else begin
          pht_1_193 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_194 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15176) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_194 <= _pht_T_3;
        end else begin
          pht_1_194 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_195 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15179) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_195 <= _pht_T_3;
        end else begin
          pht_1_195 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_196 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15182) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_196 <= _pht_T_3;
        end else begin
          pht_1_196 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_197 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15185) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_197 <= _pht_T_3;
        end else begin
          pht_1_197 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_198 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15188) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_198 <= _pht_T_3;
        end else begin
          pht_1_198 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_199 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15191) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_199 <= _pht_T_3;
        end else begin
          pht_1_199 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_200 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15194) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_200 <= _pht_T_3;
        end else begin
          pht_1_200 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_201 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15197) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_201 <= _pht_T_3;
        end else begin
          pht_1_201 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_202 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15200) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_202 <= _pht_T_3;
        end else begin
          pht_1_202 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_203 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15203) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_203 <= _pht_T_3;
        end else begin
          pht_1_203 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_204 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15206) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_204 <= _pht_T_3;
        end else begin
          pht_1_204 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_205 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15209) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_205 <= _pht_T_3;
        end else begin
          pht_1_205 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_206 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15212) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_206 <= _pht_T_3;
        end else begin
          pht_1_206 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_207 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15215) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_207 <= _pht_T_3;
        end else begin
          pht_1_207 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_208 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15218) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_208 <= _pht_T_3;
        end else begin
          pht_1_208 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_209 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15221) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_209 <= _pht_T_3;
        end else begin
          pht_1_209 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_210 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15224) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_210 <= _pht_T_3;
        end else begin
          pht_1_210 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_211 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15227) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_211 <= _pht_T_3;
        end else begin
          pht_1_211 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_212 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15230) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_212 <= _pht_T_3;
        end else begin
          pht_1_212 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_213 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15233) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_213 <= _pht_T_3;
        end else begin
          pht_1_213 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_214 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15236) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_214 <= _pht_T_3;
        end else begin
          pht_1_214 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_215 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15239) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_215 <= _pht_T_3;
        end else begin
          pht_1_215 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_216 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15242) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_216 <= _pht_T_3;
        end else begin
          pht_1_216 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_217 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15245) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_217 <= _pht_T_3;
        end else begin
          pht_1_217 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_218 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15248) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_218 <= _pht_T_3;
        end else begin
          pht_1_218 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_219 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15251) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_219 <= _pht_T_3;
        end else begin
          pht_1_219 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_220 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15254) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_220 <= _pht_T_3;
        end else begin
          pht_1_220 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_221 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15257) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_221 <= _pht_T_3;
        end else begin
          pht_1_221 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_222 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15260) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_222 <= _pht_T_3;
        end else begin
          pht_1_222 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_223 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15263) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_223 <= _pht_T_3;
        end else begin
          pht_1_223 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_224 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15266) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_224 <= _pht_T_3;
        end else begin
          pht_1_224 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_225 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15269) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_225 <= _pht_T_3;
        end else begin
          pht_1_225 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_226 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15272) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_226 <= _pht_T_3;
        end else begin
          pht_1_226 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_227 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15275) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_227 <= _pht_T_3;
        end else begin
          pht_1_227 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_228 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15278) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_228 <= _pht_T_3;
        end else begin
          pht_1_228 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_229 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15281) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_229 <= _pht_T_3;
        end else begin
          pht_1_229 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_230 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15284) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_230 <= _pht_T_3;
        end else begin
          pht_1_230 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_231 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15287) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_231 <= _pht_T_3;
        end else begin
          pht_1_231 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_232 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15290) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_232 <= _pht_T_3;
        end else begin
          pht_1_232 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_233 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15293) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_233 <= _pht_T_3;
        end else begin
          pht_1_233 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_234 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15296) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_234 <= _pht_T_3;
        end else begin
          pht_1_234 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_235 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15299) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_235 <= _pht_T_3;
        end else begin
          pht_1_235 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_236 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15302) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_236 <= _pht_T_3;
        end else begin
          pht_1_236 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_237 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15305) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_237 <= _pht_T_3;
        end else begin
          pht_1_237 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_238 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15308) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_238 <= _pht_T_3;
        end else begin
          pht_1_238 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_239 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15311) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_239 <= _pht_T_3;
        end else begin
          pht_1_239 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_240 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15314) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_240 <= _pht_T_3;
        end else begin
          pht_1_240 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_241 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15317) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_241 <= _pht_T_3;
        end else begin
          pht_1_241 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_242 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15320) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_242 <= _pht_T_3;
        end else begin
          pht_1_242 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_243 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15323) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_243 <= _pht_T_3;
        end else begin
          pht_1_243 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_244 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15326) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_244 <= _pht_T_3;
        end else begin
          pht_1_244 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_245 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15329) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_245 <= _pht_T_3;
        end else begin
          pht_1_245 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_246 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15332) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_246 <= _pht_T_3;
        end else begin
          pht_1_246 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_247 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15335) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_247 <= _pht_T_3;
        end else begin
          pht_1_247 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_248 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15338) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_248 <= _pht_T_3;
        end else begin
          pht_1_248 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_249 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15341) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_249 <= _pht_T_3;
        end else begin
          pht_1_249 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_250 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15344) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_250 <= _pht_T_3;
        end else begin
          pht_1_250 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_251 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15347) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_251 <= _pht_T_3;
        end else begin
          pht_1_251 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_252 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15350) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_252 <= _pht_T_3;
        end else begin
          pht_1_252 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_253 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15353) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_253 <= _pht_T_3;
        end else begin
          pht_1_253 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_254 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15356) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_254 <= _pht_T_3;
        end else begin
          pht_1_254 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_1_255 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_15360 & _GEN_15359) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_1_255 <= _pht_T_3;
        end else begin
          pht_1_255 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_0 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15361) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_0 <= _pht_T_3;
        end else begin
          pht_2_0 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_1 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14659) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_1 <= _pht_T_3;
        end else begin
          pht_2_1 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_2 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14661) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_2 <= _pht_T_3;
        end else begin
          pht_2_2 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_3 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14663) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_3 <= _pht_T_3;
        end else begin
          pht_2_3 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_4 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14665) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_4 <= _pht_T_3;
        end else begin
          pht_2_4 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_5 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14667) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_5 <= _pht_T_3;
        end else begin
          pht_2_5 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_6 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14669) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_6 <= _pht_T_3;
        end else begin
          pht_2_6 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_7 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14671) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_7 <= _pht_T_3;
        end else begin
          pht_2_7 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_8 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14673) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_8 <= _pht_T_3;
        end else begin
          pht_2_8 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_9 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14675) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_9 <= _pht_T_3;
        end else begin
          pht_2_9 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_10 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14677) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_10 <= _pht_T_3;
        end else begin
          pht_2_10 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_11 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14679) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_11 <= _pht_T_3;
        end else begin
          pht_2_11 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_12 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14681) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_12 <= _pht_T_3;
        end else begin
          pht_2_12 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_13 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14683) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_13 <= _pht_T_3;
        end else begin
          pht_2_13 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_14 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14685) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_14 <= _pht_T_3;
        end else begin
          pht_2_14 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_15 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14687) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_15 <= _pht_T_3;
        end else begin
          pht_2_15 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_16 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14689) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_16 <= _pht_T_3;
        end else begin
          pht_2_16 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_17 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14691) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_17 <= _pht_T_3;
        end else begin
          pht_2_17 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_18 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14693) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_18 <= _pht_T_3;
        end else begin
          pht_2_18 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_19 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14695) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_19 <= _pht_T_3;
        end else begin
          pht_2_19 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_20 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14697) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_20 <= _pht_T_3;
        end else begin
          pht_2_20 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_21 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14699) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_21 <= _pht_T_3;
        end else begin
          pht_2_21 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_22 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14701) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_22 <= _pht_T_3;
        end else begin
          pht_2_22 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_23 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14703) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_23 <= _pht_T_3;
        end else begin
          pht_2_23 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_24 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14705) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_24 <= _pht_T_3;
        end else begin
          pht_2_24 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_25 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14707) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_25 <= _pht_T_3;
        end else begin
          pht_2_25 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_26 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14709) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_26 <= _pht_T_3;
        end else begin
          pht_2_26 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_27 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14711) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_27 <= _pht_T_3;
        end else begin
          pht_2_27 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_28 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14713) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_28 <= _pht_T_3;
        end else begin
          pht_2_28 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_29 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14715) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_29 <= _pht_T_3;
        end else begin
          pht_2_29 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_30 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14717) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_30 <= _pht_T_3;
        end else begin
          pht_2_30 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_31 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14719) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_31 <= _pht_T_3;
        end else begin
          pht_2_31 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_32 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14721) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_32 <= _pht_T_3;
        end else begin
          pht_2_32 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_33 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14723) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_33 <= _pht_T_3;
        end else begin
          pht_2_33 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_34 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14725) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_34 <= _pht_T_3;
        end else begin
          pht_2_34 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_35 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14727) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_35 <= _pht_T_3;
        end else begin
          pht_2_35 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_36 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14729) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_36 <= _pht_T_3;
        end else begin
          pht_2_36 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_37 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14731) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_37 <= _pht_T_3;
        end else begin
          pht_2_37 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_38 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14733) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_38 <= _pht_T_3;
        end else begin
          pht_2_38 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_39 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14735) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_39 <= _pht_T_3;
        end else begin
          pht_2_39 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_40 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14737) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_40 <= _pht_T_3;
        end else begin
          pht_2_40 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_41 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14739) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_41 <= _pht_T_3;
        end else begin
          pht_2_41 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_42 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14741) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_42 <= _pht_T_3;
        end else begin
          pht_2_42 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_43 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14743) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_43 <= _pht_T_3;
        end else begin
          pht_2_43 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_44 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14745) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_44 <= _pht_T_3;
        end else begin
          pht_2_44 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_45 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14747) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_45 <= _pht_T_3;
        end else begin
          pht_2_45 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_46 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14749) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_46 <= _pht_T_3;
        end else begin
          pht_2_46 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_47 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14751) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_47 <= _pht_T_3;
        end else begin
          pht_2_47 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_48 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14753) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_48 <= _pht_T_3;
        end else begin
          pht_2_48 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_49 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14755) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_49 <= _pht_T_3;
        end else begin
          pht_2_49 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_50 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14757) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_50 <= _pht_T_3;
        end else begin
          pht_2_50 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_51 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14759) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_51 <= _pht_T_3;
        end else begin
          pht_2_51 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_52 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14761) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_52 <= _pht_T_3;
        end else begin
          pht_2_52 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_53 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14763) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_53 <= _pht_T_3;
        end else begin
          pht_2_53 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_54 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14765) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_54 <= _pht_T_3;
        end else begin
          pht_2_54 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_55 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14767) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_55 <= _pht_T_3;
        end else begin
          pht_2_55 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_56 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14769) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_56 <= _pht_T_3;
        end else begin
          pht_2_56 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_57 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14771) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_57 <= _pht_T_3;
        end else begin
          pht_2_57 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_58 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14773) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_58 <= _pht_T_3;
        end else begin
          pht_2_58 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_59 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14775) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_59 <= _pht_T_3;
        end else begin
          pht_2_59 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_60 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14777) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_60 <= _pht_T_3;
        end else begin
          pht_2_60 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_61 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14779) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_61 <= _pht_T_3;
        end else begin
          pht_2_61 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_62 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14781) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_62 <= _pht_T_3;
        end else begin
          pht_2_62 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_63 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14783) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_63 <= _pht_T_3;
        end else begin
          pht_2_63 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_64 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14786) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_64 <= _pht_T_3;
        end else begin
          pht_2_64 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_65 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14789) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_65 <= _pht_T_3;
        end else begin
          pht_2_65 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_66 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14792) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_66 <= _pht_T_3;
        end else begin
          pht_2_66 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_67 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14795) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_67 <= _pht_T_3;
        end else begin
          pht_2_67 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_68 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14798) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_68 <= _pht_T_3;
        end else begin
          pht_2_68 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_69 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14801) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_69 <= _pht_T_3;
        end else begin
          pht_2_69 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_70 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14804) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_70 <= _pht_T_3;
        end else begin
          pht_2_70 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_71 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14807) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_71 <= _pht_T_3;
        end else begin
          pht_2_71 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_72 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14810) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_72 <= _pht_T_3;
        end else begin
          pht_2_72 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_73 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14813) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_73 <= _pht_T_3;
        end else begin
          pht_2_73 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_74 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14816) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_74 <= _pht_T_3;
        end else begin
          pht_2_74 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_75 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14819) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_75 <= _pht_T_3;
        end else begin
          pht_2_75 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_76 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14822) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_76 <= _pht_T_3;
        end else begin
          pht_2_76 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_77 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14825) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_77 <= _pht_T_3;
        end else begin
          pht_2_77 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_78 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14828) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_78 <= _pht_T_3;
        end else begin
          pht_2_78 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_79 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14831) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_79 <= _pht_T_3;
        end else begin
          pht_2_79 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_80 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14834) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_80 <= _pht_T_3;
        end else begin
          pht_2_80 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_81 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14837) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_81 <= _pht_T_3;
        end else begin
          pht_2_81 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_82 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14840) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_82 <= _pht_T_3;
        end else begin
          pht_2_82 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_83 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14843) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_83 <= _pht_T_3;
        end else begin
          pht_2_83 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_84 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14846) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_84 <= _pht_T_3;
        end else begin
          pht_2_84 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_85 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14849) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_85 <= _pht_T_3;
        end else begin
          pht_2_85 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_86 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14852) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_86 <= _pht_T_3;
        end else begin
          pht_2_86 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_87 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14855) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_87 <= _pht_T_3;
        end else begin
          pht_2_87 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_88 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14858) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_88 <= _pht_T_3;
        end else begin
          pht_2_88 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_89 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14861) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_89 <= _pht_T_3;
        end else begin
          pht_2_89 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_90 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14864) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_90 <= _pht_T_3;
        end else begin
          pht_2_90 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_91 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14867) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_91 <= _pht_T_3;
        end else begin
          pht_2_91 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_92 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14870) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_92 <= _pht_T_3;
        end else begin
          pht_2_92 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_93 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14873) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_93 <= _pht_T_3;
        end else begin
          pht_2_93 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_94 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14876) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_94 <= _pht_T_3;
        end else begin
          pht_2_94 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_95 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14879) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_95 <= _pht_T_3;
        end else begin
          pht_2_95 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_96 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14882) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_96 <= _pht_T_3;
        end else begin
          pht_2_96 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_97 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14885) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_97 <= _pht_T_3;
        end else begin
          pht_2_97 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_98 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14888) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_98 <= _pht_T_3;
        end else begin
          pht_2_98 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_99 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14891) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_99 <= _pht_T_3;
        end else begin
          pht_2_99 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_100 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14894) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_100 <= _pht_T_3;
        end else begin
          pht_2_100 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_101 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14897) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_101 <= _pht_T_3;
        end else begin
          pht_2_101 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_102 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14900) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_102 <= _pht_T_3;
        end else begin
          pht_2_102 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_103 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14903) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_103 <= _pht_T_3;
        end else begin
          pht_2_103 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_104 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14906) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_104 <= _pht_T_3;
        end else begin
          pht_2_104 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_105 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14909) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_105 <= _pht_T_3;
        end else begin
          pht_2_105 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_106 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14912) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_106 <= _pht_T_3;
        end else begin
          pht_2_106 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_107 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14915) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_107 <= _pht_T_3;
        end else begin
          pht_2_107 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_108 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14918) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_108 <= _pht_T_3;
        end else begin
          pht_2_108 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_109 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14921) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_109 <= _pht_T_3;
        end else begin
          pht_2_109 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_110 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14924) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_110 <= _pht_T_3;
        end else begin
          pht_2_110 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_111 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14927) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_111 <= _pht_T_3;
        end else begin
          pht_2_111 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_112 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14930) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_112 <= _pht_T_3;
        end else begin
          pht_2_112 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_113 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14933) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_113 <= _pht_T_3;
        end else begin
          pht_2_113 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_114 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14936) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_114 <= _pht_T_3;
        end else begin
          pht_2_114 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_115 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14939) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_115 <= _pht_T_3;
        end else begin
          pht_2_115 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_116 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14942) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_116 <= _pht_T_3;
        end else begin
          pht_2_116 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_117 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14945) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_117 <= _pht_T_3;
        end else begin
          pht_2_117 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_118 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14948) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_118 <= _pht_T_3;
        end else begin
          pht_2_118 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_119 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14951) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_119 <= _pht_T_3;
        end else begin
          pht_2_119 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_120 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14954) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_120 <= _pht_T_3;
        end else begin
          pht_2_120 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_121 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14957) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_121 <= _pht_T_3;
        end else begin
          pht_2_121 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_122 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14960) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_122 <= _pht_T_3;
        end else begin
          pht_2_122 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_123 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14963) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_123 <= _pht_T_3;
        end else begin
          pht_2_123 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_124 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14966) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_124 <= _pht_T_3;
        end else begin
          pht_2_124 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_125 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14969) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_125 <= _pht_T_3;
        end else begin
          pht_2_125 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_126 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14972) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_126 <= _pht_T_3;
        end else begin
          pht_2_126 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_127 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14975) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_127 <= _pht_T_3;
        end else begin
          pht_2_127 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_128 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14978) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_128 <= _pht_T_3;
        end else begin
          pht_2_128 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_129 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14981) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_129 <= _pht_T_3;
        end else begin
          pht_2_129 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_130 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14984) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_130 <= _pht_T_3;
        end else begin
          pht_2_130 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_131 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14987) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_131 <= _pht_T_3;
        end else begin
          pht_2_131 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_132 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14990) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_132 <= _pht_T_3;
        end else begin
          pht_2_132 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_133 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14993) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_133 <= _pht_T_3;
        end else begin
          pht_2_133 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_134 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14996) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_134 <= _pht_T_3;
        end else begin
          pht_2_134 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_135 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_14999) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_135 <= _pht_T_3;
        end else begin
          pht_2_135 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_136 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15002) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_136 <= _pht_T_3;
        end else begin
          pht_2_136 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_137 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15005) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_137 <= _pht_T_3;
        end else begin
          pht_2_137 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_138 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15008) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_138 <= _pht_T_3;
        end else begin
          pht_2_138 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_139 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15011) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_139 <= _pht_T_3;
        end else begin
          pht_2_139 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_140 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15014) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_140 <= _pht_T_3;
        end else begin
          pht_2_140 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_141 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15017) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_141 <= _pht_T_3;
        end else begin
          pht_2_141 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_142 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15020) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_142 <= _pht_T_3;
        end else begin
          pht_2_142 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_143 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15023) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_143 <= _pht_T_3;
        end else begin
          pht_2_143 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_144 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15026) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_144 <= _pht_T_3;
        end else begin
          pht_2_144 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_145 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15029) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_145 <= _pht_T_3;
        end else begin
          pht_2_145 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_146 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15032) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_146 <= _pht_T_3;
        end else begin
          pht_2_146 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_147 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15035) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_147 <= _pht_T_3;
        end else begin
          pht_2_147 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_148 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15038) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_148 <= _pht_T_3;
        end else begin
          pht_2_148 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_149 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15041) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_149 <= _pht_T_3;
        end else begin
          pht_2_149 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_150 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15044) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_150 <= _pht_T_3;
        end else begin
          pht_2_150 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_151 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15047) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_151 <= _pht_T_3;
        end else begin
          pht_2_151 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_152 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15050) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_152 <= _pht_T_3;
        end else begin
          pht_2_152 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_153 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15053) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_153 <= _pht_T_3;
        end else begin
          pht_2_153 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_154 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15056) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_154 <= _pht_T_3;
        end else begin
          pht_2_154 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_155 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15059) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_155 <= _pht_T_3;
        end else begin
          pht_2_155 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_156 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15062) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_156 <= _pht_T_3;
        end else begin
          pht_2_156 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_157 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15065) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_157 <= _pht_T_3;
        end else begin
          pht_2_157 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_158 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15068) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_158 <= _pht_T_3;
        end else begin
          pht_2_158 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_159 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15071) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_159 <= _pht_T_3;
        end else begin
          pht_2_159 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_160 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15074) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_160 <= _pht_T_3;
        end else begin
          pht_2_160 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_161 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15077) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_161 <= _pht_T_3;
        end else begin
          pht_2_161 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_162 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15080) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_162 <= _pht_T_3;
        end else begin
          pht_2_162 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_163 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15083) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_163 <= _pht_T_3;
        end else begin
          pht_2_163 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_164 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15086) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_164 <= _pht_T_3;
        end else begin
          pht_2_164 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_165 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15089) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_165 <= _pht_T_3;
        end else begin
          pht_2_165 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_166 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15092) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_166 <= _pht_T_3;
        end else begin
          pht_2_166 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_167 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15095) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_167 <= _pht_T_3;
        end else begin
          pht_2_167 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_168 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15098) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_168 <= _pht_T_3;
        end else begin
          pht_2_168 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_169 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15101) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_169 <= _pht_T_3;
        end else begin
          pht_2_169 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_170 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15104) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_170 <= _pht_T_3;
        end else begin
          pht_2_170 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_171 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15107) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_171 <= _pht_T_3;
        end else begin
          pht_2_171 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_172 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15110) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_172 <= _pht_T_3;
        end else begin
          pht_2_172 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_173 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15113) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_173 <= _pht_T_3;
        end else begin
          pht_2_173 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_174 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15116) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_174 <= _pht_T_3;
        end else begin
          pht_2_174 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_175 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15119) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_175 <= _pht_T_3;
        end else begin
          pht_2_175 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_176 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15122) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_176 <= _pht_T_3;
        end else begin
          pht_2_176 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_177 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15125) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_177 <= _pht_T_3;
        end else begin
          pht_2_177 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_178 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15128) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_178 <= _pht_T_3;
        end else begin
          pht_2_178 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_179 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15131) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_179 <= _pht_T_3;
        end else begin
          pht_2_179 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_180 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15134) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_180 <= _pht_T_3;
        end else begin
          pht_2_180 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_181 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15137) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_181 <= _pht_T_3;
        end else begin
          pht_2_181 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_182 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15140) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_182 <= _pht_T_3;
        end else begin
          pht_2_182 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_183 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15143) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_183 <= _pht_T_3;
        end else begin
          pht_2_183 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_184 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15146) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_184 <= _pht_T_3;
        end else begin
          pht_2_184 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_185 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15149) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_185 <= _pht_T_3;
        end else begin
          pht_2_185 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_186 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15152) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_186 <= _pht_T_3;
        end else begin
          pht_2_186 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_187 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15155) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_187 <= _pht_T_3;
        end else begin
          pht_2_187 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_188 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15158) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_188 <= _pht_T_3;
        end else begin
          pht_2_188 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_189 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15161) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_189 <= _pht_T_3;
        end else begin
          pht_2_189 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_190 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15164) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_190 <= _pht_T_3;
        end else begin
          pht_2_190 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_191 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15167) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_191 <= _pht_T_3;
        end else begin
          pht_2_191 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_192 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15170) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_192 <= _pht_T_3;
        end else begin
          pht_2_192 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_193 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15173) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_193 <= _pht_T_3;
        end else begin
          pht_2_193 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_194 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15176) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_194 <= _pht_T_3;
        end else begin
          pht_2_194 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_195 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15179) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_195 <= _pht_T_3;
        end else begin
          pht_2_195 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_196 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15182) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_196 <= _pht_T_3;
        end else begin
          pht_2_196 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_197 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15185) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_197 <= _pht_T_3;
        end else begin
          pht_2_197 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_198 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15188) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_198 <= _pht_T_3;
        end else begin
          pht_2_198 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_199 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15191) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_199 <= _pht_T_3;
        end else begin
          pht_2_199 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_200 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15194) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_200 <= _pht_T_3;
        end else begin
          pht_2_200 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_201 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15197) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_201 <= _pht_T_3;
        end else begin
          pht_2_201 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_202 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15200) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_202 <= _pht_T_3;
        end else begin
          pht_2_202 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_203 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15203) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_203 <= _pht_T_3;
        end else begin
          pht_2_203 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_204 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15206) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_204 <= _pht_T_3;
        end else begin
          pht_2_204 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_205 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15209) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_205 <= _pht_T_3;
        end else begin
          pht_2_205 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_206 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15212) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_206 <= _pht_T_3;
        end else begin
          pht_2_206 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_207 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15215) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_207 <= _pht_T_3;
        end else begin
          pht_2_207 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_208 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15218) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_208 <= _pht_T_3;
        end else begin
          pht_2_208 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_209 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15221) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_209 <= _pht_T_3;
        end else begin
          pht_2_209 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_210 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15224) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_210 <= _pht_T_3;
        end else begin
          pht_2_210 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_211 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15227) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_211 <= _pht_T_3;
        end else begin
          pht_2_211 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_212 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15230) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_212 <= _pht_T_3;
        end else begin
          pht_2_212 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_213 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15233) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_213 <= _pht_T_3;
        end else begin
          pht_2_213 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_214 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15236) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_214 <= _pht_T_3;
        end else begin
          pht_2_214 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_215 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15239) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_215 <= _pht_T_3;
        end else begin
          pht_2_215 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_216 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15242) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_216 <= _pht_T_3;
        end else begin
          pht_2_216 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_217 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15245) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_217 <= _pht_T_3;
        end else begin
          pht_2_217 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_218 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15248) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_218 <= _pht_T_3;
        end else begin
          pht_2_218 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_219 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15251) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_219 <= _pht_T_3;
        end else begin
          pht_2_219 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_220 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15254) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_220 <= _pht_T_3;
        end else begin
          pht_2_220 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_221 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15257) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_221 <= _pht_T_3;
        end else begin
          pht_2_221 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_222 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15260) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_222 <= _pht_T_3;
        end else begin
          pht_2_222 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_223 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15263) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_223 <= _pht_T_3;
        end else begin
          pht_2_223 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_224 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15266) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_224 <= _pht_T_3;
        end else begin
          pht_2_224 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_225 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15269) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_225 <= _pht_T_3;
        end else begin
          pht_2_225 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_226 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15272) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_226 <= _pht_T_3;
        end else begin
          pht_2_226 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_227 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15275) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_227 <= _pht_T_3;
        end else begin
          pht_2_227 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_228 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15278) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_228 <= _pht_T_3;
        end else begin
          pht_2_228 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_229 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15281) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_229 <= _pht_T_3;
        end else begin
          pht_2_229 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_230 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15284) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_230 <= _pht_T_3;
        end else begin
          pht_2_230 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_231 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15287) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_231 <= _pht_T_3;
        end else begin
          pht_2_231 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_232 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15290) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_232 <= _pht_T_3;
        end else begin
          pht_2_232 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_233 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15293) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_233 <= _pht_T_3;
        end else begin
          pht_2_233 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_234 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15296) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_234 <= _pht_T_3;
        end else begin
          pht_2_234 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_235 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15299) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_235 <= _pht_T_3;
        end else begin
          pht_2_235 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_236 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15302) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_236 <= _pht_T_3;
        end else begin
          pht_2_236 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_237 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15305) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_237 <= _pht_T_3;
        end else begin
          pht_2_237 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_238 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15308) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_238 <= _pht_T_3;
        end else begin
          pht_2_238 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_239 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15311) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_239 <= _pht_T_3;
        end else begin
          pht_2_239 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_240 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15314) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_240 <= _pht_T_3;
        end else begin
          pht_2_240 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_241 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15317) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_241 <= _pht_T_3;
        end else begin
          pht_2_241 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_242 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15320) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_242 <= _pht_T_3;
        end else begin
          pht_2_242 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_243 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15323) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_243 <= _pht_T_3;
        end else begin
          pht_2_243 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_244 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15326) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_244 <= _pht_T_3;
        end else begin
          pht_2_244 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_245 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15329) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_245 <= _pht_T_3;
        end else begin
          pht_2_245 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_246 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15332) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_246 <= _pht_T_3;
        end else begin
          pht_2_246 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_247 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15335) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_247 <= _pht_T_3;
        end else begin
          pht_2_247 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_248 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15338) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_248 <= _pht_T_3;
        end else begin
          pht_2_248 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_249 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15341) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_249 <= _pht_T_3;
        end else begin
          pht_2_249 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_250 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15344) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_250 <= _pht_T_3;
        end else begin
          pht_2_250 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_251 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15347) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_251 <= _pht_T_3;
        end else begin
          pht_2_251 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_252 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15350) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_252 <= _pht_T_3;
        end else begin
          pht_2_252 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_253 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15353) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_253 <= _pht_T_3;
        end else begin
          pht_2_253 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_254 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15356) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_254 <= _pht_T_3;
        end else begin
          pht_2_254 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_2_255 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16064 & _GEN_15359) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_2_255 <= _pht_T_3;
        end else begin
          pht_2_255 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_0 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15361) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_0 <= _pht_T_3;
        end else begin
          pht_3_0 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_1 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14659) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_1 <= _pht_T_3;
        end else begin
          pht_3_1 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_2 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14661) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_2 <= _pht_T_3;
        end else begin
          pht_3_2 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_3 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14663) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_3 <= _pht_T_3;
        end else begin
          pht_3_3 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_4 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14665) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_4 <= _pht_T_3;
        end else begin
          pht_3_4 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_5 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14667) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_5 <= _pht_T_3;
        end else begin
          pht_3_5 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_6 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14669) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_6 <= _pht_T_3;
        end else begin
          pht_3_6 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_7 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14671) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_7 <= _pht_T_3;
        end else begin
          pht_3_7 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_8 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14673) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_8 <= _pht_T_3;
        end else begin
          pht_3_8 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_9 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14675) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_9 <= _pht_T_3;
        end else begin
          pht_3_9 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_10 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14677) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_10 <= _pht_T_3;
        end else begin
          pht_3_10 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_11 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14679) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_11 <= _pht_T_3;
        end else begin
          pht_3_11 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_12 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14681) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_12 <= _pht_T_3;
        end else begin
          pht_3_12 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_13 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14683) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_13 <= _pht_T_3;
        end else begin
          pht_3_13 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_14 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14685) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_14 <= _pht_T_3;
        end else begin
          pht_3_14 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_15 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14687) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_15 <= _pht_T_3;
        end else begin
          pht_3_15 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_16 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14689) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_16 <= _pht_T_3;
        end else begin
          pht_3_16 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_17 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14691) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_17 <= _pht_T_3;
        end else begin
          pht_3_17 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_18 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14693) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_18 <= _pht_T_3;
        end else begin
          pht_3_18 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_19 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14695) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_19 <= _pht_T_3;
        end else begin
          pht_3_19 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_20 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14697) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_20 <= _pht_T_3;
        end else begin
          pht_3_20 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_21 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14699) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_21 <= _pht_T_3;
        end else begin
          pht_3_21 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_22 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14701) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_22 <= _pht_T_3;
        end else begin
          pht_3_22 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_23 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14703) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_23 <= _pht_T_3;
        end else begin
          pht_3_23 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_24 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14705) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_24 <= _pht_T_3;
        end else begin
          pht_3_24 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_25 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14707) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_25 <= _pht_T_3;
        end else begin
          pht_3_25 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_26 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14709) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_26 <= _pht_T_3;
        end else begin
          pht_3_26 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_27 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14711) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_27 <= _pht_T_3;
        end else begin
          pht_3_27 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_28 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14713) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_28 <= _pht_T_3;
        end else begin
          pht_3_28 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_29 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14715) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_29 <= _pht_T_3;
        end else begin
          pht_3_29 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_30 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14717) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_30 <= _pht_T_3;
        end else begin
          pht_3_30 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_31 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14719) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_31 <= _pht_T_3;
        end else begin
          pht_3_31 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_32 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14721) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_32 <= _pht_T_3;
        end else begin
          pht_3_32 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_33 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14723) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_33 <= _pht_T_3;
        end else begin
          pht_3_33 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_34 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14725) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_34 <= _pht_T_3;
        end else begin
          pht_3_34 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_35 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14727) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_35 <= _pht_T_3;
        end else begin
          pht_3_35 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_36 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14729) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_36 <= _pht_T_3;
        end else begin
          pht_3_36 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_37 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14731) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_37 <= _pht_T_3;
        end else begin
          pht_3_37 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_38 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14733) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_38 <= _pht_T_3;
        end else begin
          pht_3_38 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_39 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14735) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_39 <= _pht_T_3;
        end else begin
          pht_3_39 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_40 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14737) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_40 <= _pht_T_3;
        end else begin
          pht_3_40 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_41 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14739) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_41 <= _pht_T_3;
        end else begin
          pht_3_41 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_42 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14741) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_42 <= _pht_T_3;
        end else begin
          pht_3_42 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_43 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14743) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_43 <= _pht_T_3;
        end else begin
          pht_3_43 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_44 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14745) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_44 <= _pht_T_3;
        end else begin
          pht_3_44 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_45 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14747) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_45 <= _pht_T_3;
        end else begin
          pht_3_45 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_46 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14749) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_46 <= _pht_T_3;
        end else begin
          pht_3_46 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_47 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14751) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_47 <= _pht_T_3;
        end else begin
          pht_3_47 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_48 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14753) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_48 <= _pht_T_3;
        end else begin
          pht_3_48 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_49 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14755) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_49 <= _pht_T_3;
        end else begin
          pht_3_49 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_50 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14757) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_50 <= _pht_T_3;
        end else begin
          pht_3_50 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_51 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14759) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_51 <= _pht_T_3;
        end else begin
          pht_3_51 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_52 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14761) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_52 <= _pht_T_3;
        end else begin
          pht_3_52 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_53 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14763) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_53 <= _pht_T_3;
        end else begin
          pht_3_53 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_54 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14765) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_54 <= _pht_T_3;
        end else begin
          pht_3_54 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_55 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14767) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_55 <= _pht_T_3;
        end else begin
          pht_3_55 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_56 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14769) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_56 <= _pht_T_3;
        end else begin
          pht_3_56 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_57 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14771) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_57 <= _pht_T_3;
        end else begin
          pht_3_57 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_58 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14773) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_58 <= _pht_T_3;
        end else begin
          pht_3_58 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_59 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14775) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_59 <= _pht_T_3;
        end else begin
          pht_3_59 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_60 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14777) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_60 <= _pht_T_3;
        end else begin
          pht_3_60 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_61 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14779) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_61 <= _pht_T_3;
        end else begin
          pht_3_61 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_62 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14781) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_62 <= _pht_T_3;
        end else begin
          pht_3_62 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_63 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14783) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_63 <= _pht_T_3;
        end else begin
          pht_3_63 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_64 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14786) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_64 <= _pht_T_3;
        end else begin
          pht_3_64 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_65 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14789) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_65 <= _pht_T_3;
        end else begin
          pht_3_65 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_66 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14792) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_66 <= _pht_T_3;
        end else begin
          pht_3_66 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_67 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14795) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_67 <= _pht_T_3;
        end else begin
          pht_3_67 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_68 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14798) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_68 <= _pht_T_3;
        end else begin
          pht_3_68 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_69 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14801) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_69 <= _pht_T_3;
        end else begin
          pht_3_69 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_70 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14804) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_70 <= _pht_T_3;
        end else begin
          pht_3_70 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_71 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14807) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_71 <= _pht_T_3;
        end else begin
          pht_3_71 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_72 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14810) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_72 <= _pht_T_3;
        end else begin
          pht_3_72 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_73 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14813) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_73 <= _pht_T_3;
        end else begin
          pht_3_73 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_74 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14816) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_74 <= _pht_T_3;
        end else begin
          pht_3_74 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_75 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14819) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_75 <= _pht_T_3;
        end else begin
          pht_3_75 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_76 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14822) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_76 <= _pht_T_3;
        end else begin
          pht_3_76 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_77 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14825) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_77 <= _pht_T_3;
        end else begin
          pht_3_77 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_78 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14828) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_78 <= _pht_T_3;
        end else begin
          pht_3_78 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_79 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14831) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_79 <= _pht_T_3;
        end else begin
          pht_3_79 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_80 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14834) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_80 <= _pht_T_3;
        end else begin
          pht_3_80 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_81 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14837) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_81 <= _pht_T_3;
        end else begin
          pht_3_81 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_82 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14840) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_82 <= _pht_T_3;
        end else begin
          pht_3_82 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_83 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14843) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_83 <= _pht_T_3;
        end else begin
          pht_3_83 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_84 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14846) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_84 <= _pht_T_3;
        end else begin
          pht_3_84 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_85 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14849) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_85 <= _pht_T_3;
        end else begin
          pht_3_85 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_86 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14852) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_86 <= _pht_T_3;
        end else begin
          pht_3_86 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_87 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14855) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_87 <= _pht_T_3;
        end else begin
          pht_3_87 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_88 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14858) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_88 <= _pht_T_3;
        end else begin
          pht_3_88 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_89 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14861) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_89 <= _pht_T_3;
        end else begin
          pht_3_89 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_90 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14864) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_90 <= _pht_T_3;
        end else begin
          pht_3_90 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_91 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14867) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_91 <= _pht_T_3;
        end else begin
          pht_3_91 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_92 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14870) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_92 <= _pht_T_3;
        end else begin
          pht_3_92 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_93 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14873) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_93 <= _pht_T_3;
        end else begin
          pht_3_93 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_94 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14876) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_94 <= _pht_T_3;
        end else begin
          pht_3_94 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_95 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14879) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_95 <= _pht_T_3;
        end else begin
          pht_3_95 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_96 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14882) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_96 <= _pht_T_3;
        end else begin
          pht_3_96 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_97 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14885) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_97 <= _pht_T_3;
        end else begin
          pht_3_97 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_98 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14888) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_98 <= _pht_T_3;
        end else begin
          pht_3_98 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_99 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14891) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_99 <= _pht_T_3;
        end else begin
          pht_3_99 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_100 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14894) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_100 <= _pht_T_3;
        end else begin
          pht_3_100 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_101 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14897) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_101 <= _pht_T_3;
        end else begin
          pht_3_101 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_102 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14900) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_102 <= _pht_T_3;
        end else begin
          pht_3_102 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_103 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14903) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_103 <= _pht_T_3;
        end else begin
          pht_3_103 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_104 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14906) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_104 <= _pht_T_3;
        end else begin
          pht_3_104 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_105 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14909) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_105 <= _pht_T_3;
        end else begin
          pht_3_105 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_106 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14912) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_106 <= _pht_T_3;
        end else begin
          pht_3_106 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_107 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14915) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_107 <= _pht_T_3;
        end else begin
          pht_3_107 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_108 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14918) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_108 <= _pht_T_3;
        end else begin
          pht_3_108 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_109 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14921) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_109 <= _pht_T_3;
        end else begin
          pht_3_109 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_110 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14924) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_110 <= _pht_T_3;
        end else begin
          pht_3_110 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_111 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14927) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_111 <= _pht_T_3;
        end else begin
          pht_3_111 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_112 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14930) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_112 <= _pht_T_3;
        end else begin
          pht_3_112 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_113 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14933) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_113 <= _pht_T_3;
        end else begin
          pht_3_113 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_114 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14936) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_114 <= _pht_T_3;
        end else begin
          pht_3_114 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_115 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14939) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_115 <= _pht_T_3;
        end else begin
          pht_3_115 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_116 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14942) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_116 <= _pht_T_3;
        end else begin
          pht_3_116 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_117 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14945) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_117 <= _pht_T_3;
        end else begin
          pht_3_117 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_118 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14948) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_118 <= _pht_T_3;
        end else begin
          pht_3_118 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_119 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14951) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_119 <= _pht_T_3;
        end else begin
          pht_3_119 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_120 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14954) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_120 <= _pht_T_3;
        end else begin
          pht_3_120 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_121 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14957) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_121 <= _pht_T_3;
        end else begin
          pht_3_121 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_122 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14960) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_122 <= _pht_T_3;
        end else begin
          pht_3_122 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_123 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14963) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_123 <= _pht_T_3;
        end else begin
          pht_3_123 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_124 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14966) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_124 <= _pht_T_3;
        end else begin
          pht_3_124 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_125 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14969) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_125 <= _pht_T_3;
        end else begin
          pht_3_125 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_126 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14972) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_126 <= _pht_T_3;
        end else begin
          pht_3_126 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_127 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14975) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_127 <= _pht_T_3;
        end else begin
          pht_3_127 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_128 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14978) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_128 <= _pht_T_3;
        end else begin
          pht_3_128 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_129 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14981) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_129 <= _pht_T_3;
        end else begin
          pht_3_129 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_130 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14984) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_130 <= _pht_T_3;
        end else begin
          pht_3_130 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_131 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14987) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_131 <= _pht_T_3;
        end else begin
          pht_3_131 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_132 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14990) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_132 <= _pht_T_3;
        end else begin
          pht_3_132 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_133 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14993) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_133 <= _pht_T_3;
        end else begin
          pht_3_133 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_134 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14996) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_134 <= _pht_T_3;
        end else begin
          pht_3_134 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_135 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_14999) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_135 <= _pht_T_3;
        end else begin
          pht_3_135 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_136 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15002) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_136 <= _pht_T_3;
        end else begin
          pht_3_136 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_137 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15005) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_137 <= _pht_T_3;
        end else begin
          pht_3_137 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_138 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15008) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_138 <= _pht_T_3;
        end else begin
          pht_3_138 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_139 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15011) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_139 <= _pht_T_3;
        end else begin
          pht_3_139 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_140 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15014) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_140 <= _pht_T_3;
        end else begin
          pht_3_140 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_141 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15017) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_141 <= _pht_T_3;
        end else begin
          pht_3_141 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_142 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15020) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_142 <= _pht_T_3;
        end else begin
          pht_3_142 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_143 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15023) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_143 <= _pht_T_3;
        end else begin
          pht_3_143 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_144 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15026) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_144 <= _pht_T_3;
        end else begin
          pht_3_144 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_145 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15029) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_145 <= _pht_T_3;
        end else begin
          pht_3_145 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_146 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15032) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_146 <= _pht_T_3;
        end else begin
          pht_3_146 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_147 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15035) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_147 <= _pht_T_3;
        end else begin
          pht_3_147 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_148 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15038) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_148 <= _pht_T_3;
        end else begin
          pht_3_148 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_149 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15041) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_149 <= _pht_T_3;
        end else begin
          pht_3_149 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_150 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15044) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_150 <= _pht_T_3;
        end else begin
          pht_3_150 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_151 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15047) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_151 <= _pht_T_3;
        end else begin
          pht_3_151 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_152 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15050) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_152 <= _pht_T_3;
        end else begin
          pht_3_152 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_153 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15053) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_153 <= _pht_T_3;
        end else begin
          pht_3_153 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_154 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15056) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_154 <= _pht_T_3;
        end else begin
          pht_3_154 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_155 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15059) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_155 <= _pht_T_3;
        end else begin
          pht_3_155 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_156 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15062) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_156 <= _pht_T_3;
        end else begin
          pht_3_156 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_157 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15065) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_157 <= _pht_T_3;
        end else begin
          pht_3_157 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_158 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15068) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_158 <= _pht_T_3;
        end else begin
          pht_3_158 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_159 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15071) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_159 <= _pht_T_3;
        end else begin
          pht_3_159 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_160 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15074) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_160 <= _pht_T_3;
        end else begin
          pht_3_160 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_161 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15077) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_161 <= _pht_T_3;
        end else begin
          pht_3_161 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_162 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15080) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_162 <= _pht_T_3;
        end else begin
          pht_3_162 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_163 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15083) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_163 <= _pht_T_3;
        end else begin
          pht_3_163 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_164 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15086) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_164 <= _pht_T_3;
        end else begin
          pht_3_164 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_165 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15089) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_165 <= _pht_T_3;
        end else begin
          pht_3_165 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_166 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15092) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_166 <= _pht_T_3;
        end else begin
          pht_3_166 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_167 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15095) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_167 <= _pht_T_3;
        end else begin
          pht_3_167 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_168 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15098) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_168 <= _pht_T_3;
        end else begin
          pht_3_168 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_169 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15101) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_169 <= _pht_T_3;
        end else begin
          pht_3_169 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_170 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15104) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_170 <= _pht_T_3;
        end else begin
          pht_3_170 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_171 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15107) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_171 <= _pht_T_3;
        end else begin
          pht_3_171 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_172 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15110) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_172 <= _pht_T_3;
        end else begin
          pht_3_172 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_173 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15113) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_173 <= _pht_T_3;
        end else begin
          pht_3_173 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_174 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15116) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_174 <= _pht_T_3;
        end else begin
          pht_3_174 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_175 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15119) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_175 <= _pht_T_3;
        end else begin
          pht_3_175 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_176 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15122) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_176 <= _pht_T_3;
        end else begin
          pht_3_176 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_177 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15125) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_177 <= _pht_T_3;
        end else begin
          pht_3_177 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_178 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15128) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_178 <= _pht_T_3;
        end else begin
          pht_3_178 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_179 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15131) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_179 <= _pht_T_3;
        end else begin
          pht_3_179 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_180 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15134) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_180 <= _pht_T_3;
        end else begin
          pht_3_180 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_181 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15137) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_181 <= _pht_T_3;
        end else begin
          pht_3_181 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_182 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15140) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_182 <= _pht_T_3;
        end else begin
          pht_3_182 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_183 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15143) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_183 <= _pht_T_3;
        end else begin
          pht_3_183 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_184 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15146) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_184 <= _pht_T_3;
        end else begin
          pht_3_184 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_185 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15149) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_185 <= _pht_T_3;
        end else begin
          pht_3_185 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_186 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15152) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_186 <= _pht_T_3;
        end else begin
          pht_3_186 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_187 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15155) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_187 <= _pht_T_3;
        end else begin
          pht_3_187 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_188 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15158) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_188 <= _pht_T_3;
        end else begin
          pht_3_188 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_189 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15161) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_189 <= _pht_T_3;
        end else begin
          pht_3_189 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_190 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15164) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_190 <= _pht_T_3;
        end else begin
          pht_3_190 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_191 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15167) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_191 <= _pht_T_3;
        end else begin
          pht_3_191 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_192 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15170) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_192 <= _pht_T_3;
        end else begin
          pht_3_192 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_193 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15173) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_193 <= _pht_T_3;
        end else begin
          pht_3_193 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_194 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15176) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_194 <= _pht_T_3;
        end else begin
          pht_3_194 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_195 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15179) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_195 <= _pht_T_3;
        end else begin
          pht_3_195 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_196 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15182) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_196 <= _pht_T_3;
        end else begin
          pht_3_196 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_197 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15185) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_197 <= _pht_T_3;
        end else begin
          pht_3_197 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_198 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15188) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_198 <= _pht_T_3;
        end else begin
          pht_3_198 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_199 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15191) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_199 <= _pht_T_3;
        end else begin
          pht_3_199 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_200 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15194) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_200 <= _pht_T_3;
        end else begin
          pht_3_200 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_201 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15197) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_201 <= _pht_T_3;
        end else begin
          pht_3_201 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_202 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15200) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_202 <= _pht_T_3;
        end else begin
          pht_3_202 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_203 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15203) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_203 <= _pht_T_3;
        end else begin
          pht_3_203 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_204 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15206) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_204 <= _pht_T_3;
        end else begin
          pht_3_204 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_205 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15209) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_205 <= _pht_T_3;
        end else begin
          pht_3_205 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_206 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15212) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_206 <= _pht_T_3;
        end else begin
          pht_3_206 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_207 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15215) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_207 <= _pht_T_3;
        end else begin
          pht_3_207 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_208 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15218) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_208 <= _pht_T_3;
        end else begin
          pht_3_208 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_209 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15221) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_209 <= _pht_T_3;
        end else begin
          pht_3_209 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_210 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15224) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_210 <= _pht_T_3;
        end else begin
          pht_3_210 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_211 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15227) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_211 <= _pht_T_3;
        end else begin
          pht_3_211 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_212 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15230) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_212 <= _pht_T_3;
        end else begin
          pht_3_212 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_213 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15233) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_213 <= _pht_T_3;
        end else begin
          pht_3_213 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_214 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15236) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_214 <= _pht_T_3;
        end else begin
          pht_3_214 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_215 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15239) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_215 <= _pht_T_3;
        end else begin
          pht_3_215 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_216 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15242) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_216 <= _pht_T_3;
        end else begin
          pht_3_216 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_217 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15245) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_217 <= _pht_T_3;
        end else begin
          pht_3_217 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_218 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15248) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_218 <= _pht_T_3;
        end else begin
          pht_3_218 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_219 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15251) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_219 <= _pht_T_3;
        end else begin
          pht_3_219 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_220 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15254) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_220 <= _pht_T_3;
        end else begin
          pht_3_220 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_221 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15257) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_221 <= _pht_T_3;
        end else begin
          pht_3_221 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_222 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15260) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_222 <= _pht_T_3;
        end else begin
          pht_3_222 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_223 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15263) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_223 <= _pht_T_3;
        end else begin
          pht_3_223 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_224 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15266) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_224 <= _pht_T_3;
        end else begin
          pht_3_224 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_225 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15269) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_225 <= _pht_T_3;
        end else begin
          pht_3_225 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_226 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15272) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_226 <= _pht_T_3;
        end else begin
          pht_3_226 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_227 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15275) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_227 <= _pht_T_3;
        end else begin
          pht_3_227 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_228 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15278) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_228 <= _pht_T_3;
        end else begin
          pht_3_228 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_229 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15281) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_229 <= _pht_T_3;
        end else begin
          pht_3_229 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_230 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15284) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_230 <= _pht_T_3;
        end else begin
          pht_3_230 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_231 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15287) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_231 <= _pht_T_3;
        end else begin
          pht_3_231 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_232 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15290) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_232 <= _pht_T_3;
        end else begin
          pht_3_232 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_233 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15293) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_233 <= _pht_T_3;
        end else begin
          pht_3_233 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_234 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15296) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_234 <= _pht_T_3;
        end else begin
          pht_3_234 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_235 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15299) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_235 <= _pht_T_3;
        end else begin
          pht_3_235 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_236 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15302) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_236 <= _pht_T_3;
        end else begin
          pht_3_236 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_237 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15305) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_237 <= _pht_T_3;
        end else begin
          pht_3_237 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_238 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15308) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_238 <= _pht_T_3;
        end else begin
          pht_3_238 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_239 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15311) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_239 <= _pht_T_3;
        end else begin
          pht_3_239 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_240 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15314) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_240 <= _pht_T_3;
        end else begin
          pht_3_240 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_241 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15317) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_241 <= _pht_T_3;
        end else begin
          pht_3_241 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_242 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15320) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_242 <= _pht_T_3;
        end else begin
          pht_3_242 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_243 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15323) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_243 <= _pht_T_3;
        end else begin
          pht_3_243 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_244 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15326) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_244 <= _pht_T_3;
        end else begin
          pht_3_244 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_245 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15329) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_245 <= _pht_T_3;
        end else begin
          pht_3_245 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_246 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15332) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_246 <= _pht_T_3;
        end else begin
          pht_3_246 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_247 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15335) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_247 <= _pht_T_3;
        end else begin
          pht_3_247 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_248 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15338) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_248 <= _pht_T_3;
        end else begin
          pht_3_248 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_249 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15341) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_249 <= _pht_T_3;
        end else begin
          pht_3_249 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_250 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15344) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_250 <= _pht_T_3;
        end else begin
          pht_3_250 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_251 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15347) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_251 <= _pht_T_3;
        end else begin
          pht_3_251 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_252 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15350) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_252 <= _pht_T_3;
        end else begin
          pht_3_252 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_253 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15353) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_253 <= _pht_T_3;
        end else begin
          pht_3_253 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_254 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15356) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_254 <= _pht_T_3;
        end else begin
          pht_3_254 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_3_255 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_16768 & _GEN_15359) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_3_255 <= _pht_T_3;
        end else begin
          pht_3_255 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_0 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15361) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_0 <= _pht_T_3;
        end else begin
          pht_4_0 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_1 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14659) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_1 <= _pht_T_3;
        end else begin
          pht_4_1 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_2 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14661) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_2 <= _pht_T_3;
        end else begin
          pht_4_2 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_3 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14663) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_3 <= _pht_T_3;
        end else begin
          pht_4_3 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_4 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14665) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_4 <= _pht_T_3;
        end else begin
          pht_4_4 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_5 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14667) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_5 <= _pht_T_3;
        end else begin
          pht_4_5 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_6 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14669) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_6 <= _pht_T_3;
        end else begin
          pht_4_6 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_7 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14671) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_7 <= _pht_T_3;
        end else begin
          pht_4_7 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_8 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14673) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_8 <= _pht_T_3;
        end else begin
          pht_4_8 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_9 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14675) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_9 <= _pht_T_3;
        end else begin
          pht_4_9 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_10 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14677) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_10 <= _pht_T_3;
        end else begin
          pht_4_10 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_11 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14679) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_11 <= _pht_T_3;
        end else begin
          pht_4_11 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_12 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14681) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_12 <= _pht_T_3;
        end else begin
          pht_4_12 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_13 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14683) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_13 <= _pht_T_3;
        end else begin
          pht_4_13 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_14 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14685) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_14 <= _pht_T_3;
        end else begin
          pht_4_14 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_15 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14687) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_15 <= _pht_T_3;
        end else begin
          pht_4_15 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_16 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14689) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_16 <= _pht_T_3;
        end else begin
          pht_4_16 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_17 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14691) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_17 <= _pht_T_3;
        end else begin
          pht_4_17 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_18 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14693) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_18 <= _pht_T_3;
        end else begin
          pht_4_18 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_19 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14695) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_19 <= _pht_T_3;
        end else begin
          pht_4_19 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_20 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14697) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_20 <= _pht_T_3;
        end else begin
          pht_4_20 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_21 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14699) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_21 <= _pht_T_3;
        end else begin
          pht_4_21 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_22 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14701) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_22 <= _pht_T_3;
        end else begin
          pht_4_22 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_23 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14703) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_23 <= _pht_T_3;
        end else begin
          pht_4_23 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_24 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14705) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_24 <= _pht_T_3;
        end else begin
          pht_4_24 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_25 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14707) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_25 <= _pht_T_3;
        end else begin
          pht_4_25 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_26 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14709) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_26 <= _pht_T_3;
        end else begin
          pht_4_26 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_27 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14711) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_27 <= _pht_T_3;
        end else begin
          pht_4_27 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_28 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14713) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_28 <= _pht_T_3;
        end else begin
          pht_4_28 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_29 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14715) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_29 <= _pht_T_3;
        end else begin
          pht_4_29 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_30 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14717) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_30 <= _pht_T_3;
        end else begin
          pht_4_30 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_31 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14719) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_31 <= _pht_T_3;
        end else begin
          pht_4_31 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_32 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14721) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_32 <= _pht_T_3;
        end else begin
          pht_4_32 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_33 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14723) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_33 <= _pht_T_3;
        end else begin
          pht_4_33 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_34 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14725) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_34 <= _pht_T_3;
        end else begin
          pht_4_34 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_35 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14727) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_35 <= _pht_T_3;
        end else begin
          pht_4_35 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_36 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14729) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_36 <= _pht_T_3;
        end else begin
          pht_4_36 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_37 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14731) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_37 <= _pht_T_3;
        end else begin
          pht_4_37 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_38 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14733) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_38 <= _pht_T_3;
        end else begin
          pht_4_38 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_39 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14735) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_39 <= _pht_T_3;
        end else begin
          pht_4_39 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_40 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14737) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_40 <= _pht_T_3;
        end else begin
          pht_4_40 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_41 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14739) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_41 <= _pht_T_3;
        end else begin
          pht_4_41 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_42 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14741) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_42 <= _pht_T_3;
        end else begin
          pht_4_42 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_43 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14743) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_43 <= _pht_T_3;
        end else begin
          pht_4_43 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_44 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14745) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_44 <= _pht_T_3;
        end else begin
          pht_4_44 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_45 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14747) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_45 <= _pht_T_3;
        end else begin
          pht_4_45 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_46 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14749) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_46 <= _pht_T_3;
        end else begin
          pht_4_46 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_47 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14751) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_47 <= _pht_T_3;
        end else begin
          pht_4_47 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_48 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14753) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_48 <= _pht_T_3;
        end else begin
          pht_4_48 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_49 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14755) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_49 <= _pht_T_3;
        end else begin
          pht_4_49 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_50 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14757) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_50 <= _pht_T_3;
        end else begin
          pht_4_50 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_51 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14759) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_51 <= _pht_T_3;
        end else begin
          pht_4_51 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_52 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14761) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_52 <= _pht_T_3;
        end else begin
          pht_4_52 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_53 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14763) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_53 <= _pht_T_3;
        end else begin
          pht_4_53 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_54 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14765) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_54 <= _pht_T_3;
        end else begin
          pht_4_54 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_55 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14767) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_55 <= _pht_T_3;
        end else begin
          pht_4_55 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_56 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14769) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_56 <= _pht_T_3;
        end else begin
          pht_4_56 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_57 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14771) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_57 <= _pht_T_3;
        end else begin
          pht_4_57 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_58 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14773) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_58 <= _pht_T_3;
        end else begin
          pht_4_58 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_59 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14775) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_59 <= _pht_T_3;
        end else begin
          pht_4_59 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_60 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14777) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_60 <= _pht_T_3;
        end else begin
          pht_4_60 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_61 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14779) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_61 <= _pht_T_3;
        end else begin
          pht_4_61 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_62 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14781) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_62 <= _pht_T_3;
        end else begin
          pht_4_62 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_63 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14783) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_63 <= _pht_T_3;
        end else begin
          pht_4_63 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_64 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14786) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_64 <= _pht_T_3;
        end else begin
          pht_4_64 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_65 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14789) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_65 <= _pht_T_3;
        end else begin
          pht_4_65 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_66 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14792) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_66 <= _pht_T_3;
        end else begin
          pht_4_66 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_67 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14795) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_67 <= _pht_T_3;
        end else begin
          pht_4_67 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_68 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14798) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_68 <= _pht_T_3;
        end else begin
          pht_4_68 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_69 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14801) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_69 <= _pht_T_3;
        end else begin
          pht_4_69 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_70 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14804) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_70 <= _pht_T_3;
        end else begin
          pht_4_70 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_71 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14807) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_71 <= _pht_T_3;
        end else begin
          pht_4_71 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_72 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14810) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_72 <= _pht_T_3;
        end else begin
          pht_4_72 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_73 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14813) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_73 <= _pht_T_3;
        end else begin
          pht_4_73 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_74 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14816) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_74 <= _pht_T_3;
        end else begin
          pht_4_74 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_75 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14819) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_75 <= _pht_T_3;
        end else begin
          pht_4_75 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_76 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14822) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_76 <= _pht_T_3;
        end else begin
          pht_4_76 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_77 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14825) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_77 <= _pht_T_3;
        end else begin
          pht_4_77 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_78 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14828) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_78 <= _pht_T_3;
        end else begin
          pht_4_78 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_79 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14831) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_79 <= _pht_T_3;
        end else begin
          pht_4_79 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_80 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14834) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_80 <= _pht_T_3;
        end else begin
          pht_4_80 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_81 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14837) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_81 <= _pht_T_3;
        end else begin
          pht_4_81 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_82 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14840) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_82 <= _pht_T_3;
        end else begin
          pht_4_82 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_83 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14843) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_83 <= _pht_T_3;
        end else begin
          pht_4_83 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_84 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14846) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_84 <= _pht_T_3;
        end else begin
          pht_4_84 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_85 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14849) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_85 <= _pht_T_3;
        end else begin
          pht_4_85 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_86 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14852) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_86 <= _pht_T_3;
        end else begin
          pht_4_86 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_87 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14855) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_87 <= _pht_T_3;
        end else begin
          pht_4_87 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_88 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14858) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_88 <= _pht_T_3;
        end else begin
          pht_4_88 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_89 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14861) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_89 <= _pht_T_3;
        end else begin
          pht_4_89 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_90 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14864) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_90 <= _pht_T_3;
        end else begin
          pht_4_90 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_91 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14867) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_91 <= _pht_T_3;
        end else begin
          pht_4_91 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_92 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14870) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_92 <= _pht_T_3;
        end else begin
          pht_4_92 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_93 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14873) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_93 <= _pht_T_3;
        end else begin
          pht_4_93 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_94 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14876) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_94 <= _pht_T_3;
        end else begin
          pht_4_94 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_95 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14879) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_95 <= _pht_T_3;
        end else begin
          pht_4_95 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_96 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14882) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_96 <= _pht_T_3;
        end else begin
          pht_4_96 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_97 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14885) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_97 <= _pht_T_3;
        end else begin
          pht_4_97 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_98 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14888) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_98 <= _pht_T_3;
        end else begin
          pht_4_98 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_99 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14891) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_99 <= _pht_T_3;
        end else begin
          pht_4_99 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_100 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14894) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_100 <= _pht_T_3;
        end else begin
          pht_4_100 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_101 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14897) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_101 <= _pht_T_3;
        end else begin
          pht_4_101 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_102 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14900) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_102 <= _pht_T_3;
        end else begin
          pht_4_102 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_103 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14903) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_103 <= _pht_T_3;
        end else begin
          pht_4_103 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_104 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14906) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_104 <= _pht_T_3;
        end else begin
          pht_4_104 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_105 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14909) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_105 <= _pht_T_3;
        end else begin
          pht_4_105 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_106 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14912) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_106 <= _pht_T_3;
        end else begin
          pht_4_106 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_107 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14915) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_107 <= _pht_T_3;
        end else begin
          pht_4_107 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_108 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14918) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_108 <= _pht_T_3;
        end else begin
          pht_4_108 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_109 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14921) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_109 <= _pht_T_3;
        end else begin
          pht_4_109 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_110 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14924) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_110 <= _pht_T_3;
        end else begin
          pht_4_110 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_111 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14927) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_111 <= _pht_T_3;
        end else begin
          pht_4_111 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_112 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14930) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_112 <= _pht_T_3;
        end else begin
          pht_4_112 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_113 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14933) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_113 <= _pht_T_3;
        end else begin
          pht_4_113 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_114 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14936) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_114 <= _pht_T_3;
        end else begin
          pht_4_114 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_115 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14939) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_115 <= _pht_T_3;
        end else begin
          pht_4_115 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_116 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14942) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_116 <= _pht_T_3;
        end else begin
          pht_4_116 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_117 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14945) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_117 <= _pht_T_3;
        end else begin
          pht_4_117 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_118 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14948) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_118 <= _pht_T_3;
        end else begin
          pht_4_118 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_119 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14951) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_119 <= _pht_T_3;
        end else begin
          pht_4_119 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_120 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14954) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_120 <= _pht_T_3;
        end else begin
          pht_4_120 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_121 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14957) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_121 <= _pht_T_3;
        end else begin
          pht_4_121 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_122 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14960) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_122 <= _pht_T_3;
        end else begin
          pht_4_122 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_123 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14963) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_123 <= _pht_T_3;
        end else begin
          pht_4_123 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_124 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14966) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_124 <= _pht_T_3;
        end else begin
          pht_4_124 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_125 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14969) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_125 <= _pht_T_3;
        end else begin
          pht_4_125 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_126 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14972) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_126 <= _pht_T_3;
        end else begin
          pht_4_126 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_127 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14975) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_127 <= _pht_T_3;
        end else begin
          pht_4_127 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_128 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14978) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_128 <= _pht_T_3;
        end else begin
          pht_4_128 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_129 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14981) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_129 <= _pht_T_3;
        end else begin
          pht_4_129 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_130 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14984) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_130 <= _pht_T_3;
        end else begin
          pht_4_130 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_131 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14987) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_131 <= _pht_T_3;
        end else begin
          pht_4_131 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_132 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14990) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_132 <= _pht_T_3;
        end else begin
          pht_4_132 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_133 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14993) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_133 <= _pht_T_3;
        end else begin
          pht_4_133 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_134 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14996) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_134 <= _pht_T_3;
        end else begin
          pht_4_134 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_135 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_14999) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_135 <= _pht_T_3;
        end else begin
          pht_4_135 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_136 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15002) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_136 <= _pht_T_3;
        end else begin
          pht_4_136 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_137 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15005) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_137 <= _pht_T_3;
        end else begin
          pht_4_137 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_138 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15008) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_138 <= _pht_T_3;
        end else begin
          pht_4_138 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_139 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15011) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_139 <= _pht_T_3;
        end else begin
          pht_4_139 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_140 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15014) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_140 <= _pht_T_3;
        end else begin
          pht_4_140 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_141 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15017) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_141 <= _pht_T_3;
        end else begin
          pht_4_141 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_142 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15020) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_142 <= _pht_T_3;
        end else begin
          pht_4_142 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_143 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15023) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_143 <= _pht_T_3;
        end else begin
          pht_4_143 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_144 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15026) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_144 <= _pht_T_3;
        end else begin
          pht_4_144 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_145 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15029) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_145 <= _pht_T_3;
        end else begin
          pht_4_145 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_146 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15032) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_146 <= _pht_T_3;
        end else begin
          pht_4_146 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_147 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15035) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_147 <= _pht_T_3;
        end else begin
          pht_4_147 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_148 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15038) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_148 <= _pht_T_3;
        end else begin
          pht_4_148 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_149 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15041) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_149 <= _pht_T_3;
        end else begin
          pht_4_149 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_150 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15044) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_150 <= _pht_T_3;
        end else begin
          pht_4_150 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_151 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15047) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_151 <= _pht_T_3;
        end else begin
          pht_4_151 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_152 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15050) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_152 <= _pht_T_3;
        end else begin
          pht_4_152 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_153 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15053) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_153 <= _pht_T_3;
        end else begin
          pht_4_153 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_154 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15056) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_154 <= _pht_T_3;
        end else begin
          pht_4_154 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_155 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15059) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_155 <= _pht_T_3;
        end else begin
          pht_4_155 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_156 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15062) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_156 <= _pht_T_3;
        end else begin
          pht_4_156 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_157 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15065) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_157 <= _pht_T_3;
        end else begin
          pht_4_157 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_158 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15068) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_158 <= _pht_T_3;
        end else begin
          pht_4_158 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_159 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15071) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_159 <= _pht_T_3;
        end else begin
          pht_4_159 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_160 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15074) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_160 <= _pht_T_3;
        end else begin
          pht_4_160 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_161 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15077) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_161 <= _pht_T_3;
        end else begin
          pht_4_161 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_162 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15080) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_162 <= _pht_T_3;
        end else begin
          pht_4_162 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_163 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15083) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_163 <= _pht_T_3;
        end else begin
          pht_4_163 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_164 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15086) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_164 <= _pht_T_3;
        end else begin
          pht_4_164 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_165 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15089) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_165 <= _pht_T_3;
        end else begin
          pht_4_165 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_166 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15092) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_166 <= _pht_T_3;
        end else begin
          pht_4_166 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_167 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15095) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_167 <= _pht_T_3;
        end else begin
          pht_4_167 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_168 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15098) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_168 <= _pht_T_3;
        end else begin
          pht_4_168 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_169 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15101) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_169 <= _pht_T_3;
        end else begin
          pht_4_169 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_170 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15104) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_170 <= _pht_T_3;
        end else begin
          pht_4_170 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_171 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15107) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_171 <= _pht_T_3;
        end else begin
          pht_4_171 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_172 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15110) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_172 <= _pht_T_3;
        end else begin
          pht_4_172 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_173 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15113) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_173 <= _pht_T_3;
        end else begin
          pht_4_173 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_174 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15116) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_174 <= _pht_T_3;
        end else begin
          pht_4_174 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_175 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15119) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_175 <= _pht_T_3;
        end else begin
          pht_4_175 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_176 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15122) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_176 <= _pht_T_3;
        end else begin
          pht_4_176 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_177 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15125) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_177 <= _pht_T_3;
        end else begin
          pht_4_177 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_178 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15128) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_178 <= _pht_T_3;
        end else begin
          pht_4_178 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_179 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15131) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_179 <= _pht_T_3;
        end else begin
          pht_4_179 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_180 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15134) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_180 <= _pht_T_3;
        end else begin
          pht_4_180 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_181 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15137) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_181 <= _pht_T_3;
        end else begin
          pht_4_181 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_182 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15140) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_182 <= _pht_T_3;
        end else begin
          pht_4_182 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_183 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15143) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_183 <= _pht_T_3;
        end else begin
          pht_4_183 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_184 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15146) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_184 <= _pht_T_3;
        end else begin
          pht_4_184 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_185 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15149) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_185 <= _pht_T_3;
        end else begin
          pht_4_185 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_186 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15152) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_186 <= _pht_T_3;
        end else begin
          pht_4_186 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_187 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15155) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_187 <= _pht_T_3;
        end else begin
          pht_4_187 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_188 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15158) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_188 <= _pht_T_3;
        end else begin
          pht_4_188 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_189 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15161) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_189 <= _pht_T_3;
        end else begin
          pht_4_189 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_190 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15164) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_190 <= _pht_T_3;
        end else begin
          pht_4_190 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_191 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15167) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_191 <= _pht_T_3;
        end else begin
          pht_4_191 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_192 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15170) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_192 <= _pht_T_3;
        end else begin
          pht_4_192 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_193 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15173) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_193 <= _pht_T_3;
        end else begin
          pht_4_193 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_194 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15176) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_194 <= _pht_T_3;
        end else begin
          pht_4_194 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_195 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15179) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_195 <= _pht_T_3;
        end else begin
          pht_4_195 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_196 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15182) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_196 <= _pht_T_3;
        end else begin
          pht_4_196 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_197 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15185) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_197 <= _pht_T_3;
        end else begin
          pht_4_197 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_198 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15188) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_198 <= _pht_T_3;
        end else begin
          pht_4_198 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_199 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15191) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_199 <= _pht_T_3;
        end else begin
          pht_4_199 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_200 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15194) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_200 <= _pht_T_3;
        end else begin
          pht_4_200 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_201 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15197) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_201 <= _pht_T_3;
        end else begin
          pht_4_201 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_202 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15200) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_202 <= _pht_T_3;
        end else begin
          pht_4_202 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_203 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15203) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_203 <= _pht_T_3;
        end else begin
          pht_4_203 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_204 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15206) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_204 <= _pht_T_3;
        end else begin
          pht_4_204 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_205 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15209) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_205 <= _pht_T_3;
        end else begin
          pht_4_205 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_206 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15212) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_206 <= _pht_T_3;
        end else begin
          pht_4_206 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_207 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15215) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_207 <= _pht_T_3;
        end else begin
          pht_4_207 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_208 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15218) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_208 <= _pht_T_3;
        end else begin
          pht_4_208 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_209 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15221) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_209 <= _pht_T_3;
        end else begin
          pht_4_209 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_210 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15224) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_210 <= _pht_T_3;
        end else begin
          pht_4_210 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_211 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15227) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_211 <= _pht_T_3;
        end else begin
          pht_4_211 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_212 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15230) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_212 <= _pht_T_3;
        end else begin
          pht_4_212 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_213 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15233) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_213 <= _pht_T_3;
        end else begin
          pht_4_213 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_214 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15236) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_214 <= _pht_T_3;
        end else begin
          pht_4_214 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_215 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15239) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_215 <= _pht_T_3;
        end else begin
          pht_4_215 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_216 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15242) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_216 <= _pht_T_3;
        end else begin
          pht_4_216 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_217 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15245) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_217 <= _pht_T_3;
        end else begin
          pht_4_217 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_218 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15248) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_218 <= _pht_T_3;
        end else begin
          pht_4_218 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_219 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15251) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_219 <= _pht_T_3;
        end else begin
          pht_4_219 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_220 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15254) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_220 <= _pht_T_3;
        end else begin
          pht_4_220 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_221 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15257) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_221 <= _pht_T_3;
        end else begin
          pht_4_221 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_222 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15260) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_222 <= _pht_T_3;
        end else begin
          pht_4_222 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_223 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15263) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_223 <= _pht_T_3;
        end else begin
          pht_4_223 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_224 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15266) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_224 <= _pht_T_3;
        end else begin
          pht_4_224 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_225 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15269) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_225 <= _pht_T_3;
        end else begin
          pht_4_225 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_226 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15272) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_226 <= _pht_T_3;
        end else begin
          pht_4_226 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_227 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15275) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_227 <= _pht_T_3;
        end else begin
          pht_4_227 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_228 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15278) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_228 <= _pht_T_3;
        end else begin
          pht_4_228 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_229 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15281) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_229 <= _pht_T_3;
        end else begin
          pht_4_229 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_230 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15284) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_230 <= _pht_T_3;
        end else begin
          pht_4_230 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_231 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15287) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_231 <= _pht_T_3;
        end else begin
          pht_4_231 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_232 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15290) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_232 <= _pht_T_3;
        end else begin
          pht_4_232 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_233 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15293) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_233 <= _pht_T_3;
        end else begin
          pht_4_233 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_234 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15296) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_234 <= _pht_T_3;
        end else begin
          pht_4_234 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_235 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15299) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_235 <= _pht_T_3;
        end else begin
          pht_4_235 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_236 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15302) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_236 <= _pht_T_3;
        end else begin
          pht_4_236 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_237 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15305) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_237 <= _pht_T_3;
        end else begin
          pht_4_237 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_238 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15308) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_238 <= _pht_T_3;
        end else begin
          pht_4_238 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_239 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15311) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_239 <= _pht_T_3;
        end else begin
          pht_4_239 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_240 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15314) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_240 <= _pht_T_3;
        end else begin
          pht_4_240 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_241 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15317) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_241 <= _pht_T_3;
        end else begin
          pht_4_241 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_242 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15320) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_242 <= _pht_T_3;
        end else begin
          pht_4_242 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_243 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15323) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_243 <= _pht_T_3;
        end else begin
          pht_4_243 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_244 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15326) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_244 <= _pht_T_3;
        end else begin
          pht_4_244 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_245 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15329) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_245 <= _pht_T_3;
        end else begin
          pht_4_245 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_246 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15332) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_246 <= _pht_T_3;
        end else begin
          pht_4_246 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_247 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15335) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_247 <= _pht_T_3;
        end else begin
          pht_4_247 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_248 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15338) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_248 <= _pht_T_3;
        end else begin
          pht_4_248 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_249 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15341) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_249 <= _pht_T_3;
        end else begin
          pht_4_249 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_250 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15344) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_250 <= _pht_T_3;
        end else begin
          pht_4_250 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_251 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15347) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_251 <= _pht_T_3;
        end else begin
          pht_4_251 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_252 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15350) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_252 <= _pht_T_3;
        end else begin
          pht_4_252 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_253 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15353) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_253 <= _pht_T_3;
        end else begin
          pht_4_253 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_254 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15356) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_254 <= _pht_T_3;
        end else begin
          pht_4_254 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_4_255 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_17472 & _GEN_15359) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_4_255 <= _pht_T_3;
        end else begin
          pht_4_255 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_0 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15361) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_0 <= _pht_T_3;
        end else begin
          pht_5_0 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_1 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14659) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_1 <= _pht_T_3;
        end else begin
          pht_5_1 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_2 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14661) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_2 <= _pht_T_3;
        end else begin
          pht_5_2 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_3 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14663) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_3 <= _pht_T_3;
        end else begin
          pht_5_3 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_4 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14665) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_4 <= _pht_T_3;
        end else begin
          pht_5_4 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_5 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14667) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_5 <= _pht_T_3;
        end else begin
          pht_5_5 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_6 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14669) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_6 <= _pht_T_3;
        end else begin
          pht_5_6 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_7 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14671) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_7 <= _pht_T_3;
        end else begin
          pht_5_7 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_8 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14673) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_8 <= _pht_T_3;
        end else begin
          pht_5_8 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_9 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14675) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_9 <= _pht_T_3;
        end else begin
          pht_5_9 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_10 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14677) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_10 <= _pht_T_3;
        end else begin
          pht_5_10 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_11 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14679) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_11 <= _pht_T_3;
        end else begin
          pht_5_11 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_12 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14681) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_12 <= _pht_T_3;
        end else begin
          pht_5_12 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_13 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14683) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_13 <= _pht_T_3;
        end else begin
          pht_5_13 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_14 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14685) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_14 <= _pht_T_3;
        end else begin
          pht_5_14 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_15 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14687) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_15 <= _pht_T_3;
        end else begin
          pht_5_15 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_16 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14689) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_16 <= _pht_T_3;
        end else begin
          pht_5_16 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_17 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14691) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_17 <= _pht_T_3;
        end else begin
          pht_5_17 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_18 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14693) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_18 <= _pht_T_3;
        end else begin
          pht_5_18 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_19 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14695) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_19 <= _pht_T_3;
        end else begin
          pht_5_19 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_20 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14697) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_20 <= _pht_T_3;
        end else begin
          pht_5_20 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_21 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14699) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_21 <= _pht_T_3;
        end else begin
          pht_5_21 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_22 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14701) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_22 <= _pht_T_3;
        end else begin
          pht_5_22 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_23 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14703) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_23 <= _pht_T_3;
        end else begin
          pht_5_23 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_24 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14705) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_24 <= _pht_T_3;
        end else begin
          pht_5_24 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_25 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14707) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_25 <= _pht_T_3;
        end else begin
          pht_5_25 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_26 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14709) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_26 <= _pht_T_3;
        end else begin
          pht_5_26 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_27 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14711) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_27 <= _pht_T_3;
        end else begin
          pht_5_27 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_28 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14713) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_28 <= _pht_T_3;
        end else begin
          pht_5_28 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_29 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14715) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_29 <= _pht_T_3;
        end else begin
          pht_5_29 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_30 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14717) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_30 <= _pht_T_3;
        end else begin
          pht_5_30 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_31 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14719) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_31 <= _pht_T_3;
        end else begin
          pht_5_31 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_32 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14721) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_32 <= _pht_T_3;
        end else begin
          pht_5_32 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_33 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14723) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_33 <= _pht_T_3;
        end else begin
          pht_5_33 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_34 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14725) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_34 <= _pht_T_3;
        end else begin
          pht_5_34 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_35 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14727) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_35 <= _pht_T_3;
        end else begin
          pht_5_35 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_36 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14729) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_36 <= _pht_T_3;
        end else begin
          pht_5_36 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_37 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14731) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_37 <= _pht_T_3;
        end else begin
          pht_5_37 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_38 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14733) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_38 <= _pht_T_3;
        end else begin
          pht_5_38 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_39 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14735) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_39 <= _pht_T_3;
        end else begin
          pht_5_39 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_40 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14737) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_40 <= _pht_T_3;
        end else begin
          pht_5_40 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_41 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14739) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_41 <= _pht_T_3;
        end else begin
          pht_5_41 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_42 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14741) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_42 <= _pht_T_3;
        end else begin
          pht_5_42 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_43 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14743) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_43 <= _pht_T_3;
        end else begin
          pht_5_43 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_44 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14745) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_44 <= _pht_T_3;
        end else begin
          pht_5_44 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_45 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14747) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_45 <= _pht_T_3;
        end else begin
          pht_5_45 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_46 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14749) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_46 <= _pht_T_3;
        end else begin
          pht_5_46 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_47 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14751) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_47 <= _pht_T_3;
        end else begin
          pht_5_47 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_48 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14753) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_48 <= _pht_T_3;
        end else begin
          pht_5_48 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_49 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14755) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_49 <= _pht_T_3;
        end else begin
          pht_5_49 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_50 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14757) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_50 <= _pht_T_3;
        end else begin
          pht_5_50 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_51 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14759) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_51 <= _pht_T_3;
        end else begin
          pht_5_51 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_52 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14761) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_52 <= _pht_T_3;
        end else begin
          pht_5_52 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_53 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14763) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_53 <= _pht_T_3;
        end else begin
          pht_5_53 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_54 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14765) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_54 <= _pht_T_3;
        end else begin
          pht_5_54 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_55 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14767) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_55 <= _pht_T_3;
        end else begin
          pht_5_55 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_56 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14769) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_56 <= _pht_T_3;
        end else begin
          pht_5_56 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_57 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14771) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_57 <= _pht_T_3;
        end else begin
          pht_5_57 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_58 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14773) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_58 <= _pht_T_3;
        end else begin
          pht_5_58 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_59 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14775) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_59 <= _pht_T_3;
        end else begin
          pht_5_59 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_60 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14777) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_60 <= _pht_T_3;
        end else begin
          pht_5_60 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_61 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14779) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_61 <= _pht_T_3;
        end else begin
          pht_5_61 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_62 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14781) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_62 <= _pht_T_3;
        end else begin
          pht_5_62 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_63 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14783) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_63 <= _pht_T_3;
        end else begin
          pht_5_63 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_64 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14786) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_64 <= _pht_T_3;
        end else begin
          pht_5_64 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_65 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14789) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_65 <= _pht_T_3;
        end else begin
          pht_5_65 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_66 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14792) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_66 <= _pht_T_3;
        end else begin
          pht_5_66 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_67 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14795) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_67 <= _pht_T_3;
        end else begin
          pht_5_67 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_68 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14798) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_68 <= _pht_T_3;
        end else begin
          pht_5_68 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_69 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14801) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_69 <= _pht_T_3;
        end else begin
          pht_5_69 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_70 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14804) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_70 <= _pht_T_3;
        end else begin
          pht_5_70 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_71 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14807) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_71 <= _pht_T_3;
        end else begin
          pht_5_71 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_72 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14810) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_72 <= _pht_T_3;
        end else begin
          pht_5_72 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_73 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14813) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_73 <= _pht_T_3;
        end else begin
          pht_5_73 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_74 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14816) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_74 <= _pht_T_3;
        end else begin
          pht_5_74 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_75 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14819) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_75 <= _pht_T_3;
        end else begin
          pht_5_75 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_76 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14822) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_76 <= _pht_T_3;
        end else begin
          pht_5_76 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_77 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14825) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_77 <= _pht_T_3;
        end else begin
          pht_5_77 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_78 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14828) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_78 <= _pht_T_3;
        end else begin
          pht_5_78 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_79 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14831) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_79 <= _pht_T_3;
        end else begin
          pht_5_79 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_80 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14834) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_80 <= _pht_T_3;
        end else begin
          pht_5_80 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_81 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14837) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_81 <= _pht_T_3;
        end else begin
          pht_5_81 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_82 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14840) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_82 <= _pht_T_3;
        end else begin
          pht_5_82 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_83 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14843) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_83 <= _pht_T_3;
        end else begin
          pht_5_83 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_84 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14846) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_84 <= _pht_T_3;
        end else begin
          pht_5_84 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_85 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14849) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_85 <= _pht_T_3;
        end else begin
          pht_5_85 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_86 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14852) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_86 <= _pht_T_3;
        end else begin
          pht_5_86 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_87 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14855) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_87 <= _pht_T_3;
        end else begin
          pht_5_87 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_88 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14858) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_88 <= _pht_T_3;
        end else begin
          pht_5_88 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_89 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14861) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_89 <= _pht_T_3;
        end else begin
          pht_5_89 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_90 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14864) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_90 <= _pht_T_3;
        end else begin
          pht_5_90 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_91 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14867) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_91 <= _pht_T_3;
        end else begin
          pht_5_91 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_92 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14870) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_92 <= _pht_T_3;
        end else begin
          pht_5_92 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_93 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14873) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_93 <= _pht_T_3;
        end else begin
          pht_5_93 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_94 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14876) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_94 <= _pht_T_3;
        end else begin
          pht_5_94 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_95 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14879) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_95 <= _pht_T_3;
        end else begin
          pht_5_95 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_96 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14882) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_96 <= _pht_T_3;
        end else begin
          pht_5_96 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_97 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14885) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_97 <= _pht_T_3;
        end else begin
          pht_5_97 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_98 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14888) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_98 <= _pht_T_3;
        end else begin
          pht_5_98 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_99 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14891) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_99 <= _pht_T_3;
        end else begin
          pht_5_99 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_100 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14894) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_100 <= _pht_T_3;
        end else begin
          pht_5_100 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_101 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14897) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_101 <= _pht_T_3;
        end else begin
          pht_5_101 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_102 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14900) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_102 <= _pht_T_3;
        end else begin
          pht_5_102 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_103 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14903) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_103 <= _pht_T_3;
        end else begin
          pht_5_103 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_104 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14906) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_104 <= _pht_T_3;
        end else begin
          pht_5_104 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_105 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14909) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_105 <= _pht_T_3;
        end else begin
          pht_5_105 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_106 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14912) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_106 <= _pht_T_3;
        end else begin
          pht_5_106 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_107 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14915) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_107 <= _pht_T_3;
        end else begin
          pht_5_107 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_108 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14918) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_108 <= _pht_T_3;
        end else begin
          pht_5_108 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_109 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14921) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_109 <= _pht_T_3;
        end else begin
          pht_5_109 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_110 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14924) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_110 <= _pht_T_3;
        end else begin
          pht_5_110 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_111 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14927) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_111 <= _pht_T_3;
        end else begin
          pht_5_111 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_112 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14930) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_112 <= _pht_T_3;
        end else begin
          pht_5_112 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_113 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14933) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_113 <= _pht_T_3;
        end else begin
          pht_5_113 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_114 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14936) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_114 <= _pht_T_3;
        end else begin
          pht_5_114 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_115 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14939) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_115 <= _pht_T_3;
        end else begin
          pht_5_115 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_116 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14942) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_116 <= _pht_T_3;
        end else begin
          pht_5_116 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_117 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14945) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_117 <= _pht_T_3;
        end else begin
          pht_5_117 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_118 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14948) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_118 <= _pht_T_3;
        end else begin
          pht_5_118 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_119 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14951) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_119 <= _pht_T_3;
        end else begin
          pht_5_119 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_120 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14954) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_120 <= _pht_T_3;
        end else begin
          pht_5_120 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_121 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14957) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_121 <= _pht_T_3;
        end else begin
          pht_5_121 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_122 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14960) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_122 <= _pht_T_3;
        end else begin
          pht_5_122 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_123 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14963) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_123 <= _pht_T_3;
        end else begin
          pht_5_123 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_124 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14966) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_124 <= _pht_T_3;
        end else begin
          pht_5_124 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_125 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14969) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_125 <= _pht_T_3;
        end else begin
          pht_5_125 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_126 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14972) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_126 <= _pht_T_3;
        end else begin
          pht_5_126 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_127 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14975) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_127 <= _pht_T_3;
        end else begin
          pht_5_127 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_128 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14978) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_128 <= _pht_T_3;
        end else begin
          pht_5_128 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_129 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14981) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_129 <= _pht_T_3;
        end else begin
          pht_5_129 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_130 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14984) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_130 <= _pht_T_3;
        end else begin
          pht_5_130 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_131 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14987) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_131 <= _pht_T_3;
        end else begin
          pht_5_131 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_132 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14990) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_132 <= _pht_T_3;
        end else begin
          pht_5_132 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_133 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14993) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_133 <= _pht_T_3;
        end else begin
          pht_5_133 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_134 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14996) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_134 <= _pht_T_3;
        end else begin
          pht_5_134 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_135 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_14999) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_135 <= _pht_T_3;
        end else begin
          pht_5_135 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_136 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15002) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_136 <= _pht_T_3;
        end else begin
          pht_5_136 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_137 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15005) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_137 <= _pht_T_3;
        end else begin
          pht_5_137 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_138 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15008) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_138 <= _pht_T_3;
        end else begin
          pht_5_138 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_139 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15011) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_139 <= _pht_T_3;
        end else begin
          pht_5_139 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_140 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15014) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_140 <= _pht_T_3;
        end else begin
          pht_5_140 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_141 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15017) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_141 <= _pht_T_3;
        end else begin
          pht_5_141 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_142 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15020) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_142 <= _pht_T_3;
        end else begin
          pht_5_142 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_143 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15023) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_143 <= _pht_T_3;
        end else begin
          pht_5_143 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_144 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15026) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_144 <= _pht_T_3;
        end else begin
          pht_5_144 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_145 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15029) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_145 <= _pht_T_3;
        end else begin
          pht_5_145 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_146 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15032) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_146 <= _pht_T_3;
        end else begin
          pht_5_146 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_147 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15035) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_147 <= _pht_T_3;
        end else begin
          pht_5_147 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_148 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15038) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_148 <= _pht_T_3;
        end else begin
          pht_5_148 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_149 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15041) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_149 <= _pht_T_3;
        end else begin
          pht_5_149 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_150 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15044) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_150 <= _pht_T_3;
        end else begin
          pht_5_150 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_151 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15047) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_151 <= _pht_T_3;
        end else begin
          pht_5_151 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_152 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15050) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_152 <= _pht_T_3;
        end else begin
          pht_5_152 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_153 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15053) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_153 <= _pht_T_3;
        end else begin
          pht_5_153 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_154 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15056) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_154 <= _pht_T_3;
        end else begin
          pht_5_154 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_155 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15059) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_155 <= _pht_T_3;
        end else begin
          pht_5_155 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_156 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15062) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_156 <= _pht_T_3;
        end else begin
          pht_5_156 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_157 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15065) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_157 <= _pht_T_3;
        end else begin
          pht_5_157 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_158 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15068) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_158 <= _pht_T_3;
        end else begin
          pht_5_158 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_159 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15071) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_159 <= _pht_T_3;
        end else begin
          pht_5_159 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_160 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15074) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_160 <= _pht_T_3;
        end else begin
          pht_5_160 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_161 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15077) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_161 <= _pht_T_3;
        end else begin
          pht_5_161 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_162 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15080) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_162 <= _pht_T_3;
        end else begin
          pht_5_162 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_163 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15083) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_163 <= _pht_T_3;
        end else begin
          pht_5_163 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_164 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15086) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_164 <= _pht_T_3;
        end else begin
          pht_5_164 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_165 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15089) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_165 <= _pht_T_3;
        end else begin
          pht_5_165 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_166 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15092) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_166 <= _pht_T_3;
        end else begin
          pht_5_166 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_167 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15095) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_167 <= _pht_T_3;
        end else begin
          pht_5_167 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_168 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15098) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_168 <= _pht_T_3;
        end else begin
          pht_5_168 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_169 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15101) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_169 <= _pht_T_3;
        end else begin
          pht_5_169 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_170 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15104) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_170 <= _pht_T_3;
        end else begin
          pht_5_170 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_171 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15107) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_171 <= _pht_T_3;
        end else begin
          pht_5_171 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_172 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15110) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_172 <= _pht_T_3;
        end else begin
          pht_5_172 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_173 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15113) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_173 <= _pht_T_3;
        end else begin
          pht_5_173 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_174 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15116) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_174 <= _pht_T_3;
        end else begin
          pht_5_174 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_175 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15119) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_175 <= _pht_T_3;
        end else begin
          pht_5_175 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_176 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15122) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_176 <= _pht_T_3;
        end else begin
          pht_5_176 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_177 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15125) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_177 <= _pht_T_3;
        end else begin
          pht_5_177 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_178 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15128) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_178 <= _pht_T_3;
        end else begin
          pht_5_178 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_179 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15131) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_179 <= _pht_T_3;
        end else begin
          pht_5_179 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_180 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15134) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_180 <= _pht_T_3;
        end else begin
          pht_5_180 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_181 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15137) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_181 <= _pht_T_3;
        end else begin
          pht_5_181 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_182 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15140) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_182 <= _pht_T_3;
        end else begin
          pht_5_182 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_183 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15143) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_183 <= _pht_T_3;
        end else begin
          pht_5_183 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_184 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15146) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_184 <= _pht_T_3;
        end else begin
          pht_5_184 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_185 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15149) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_185 <= _pht_T_3;
        end else begin
          pht_5_185 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_186 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15152) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_186 <= _pht_T_3;
        end else begin
          pht_5_186 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_187 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15155) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_187 <= _pht_T_3;
        end else begin
          pht_5_187 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_188 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15158) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_188 <= _pht_T_3;
        end else begin
          pht_5_188 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_189 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15161) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_189 <= _pht_T_3;
        end else begin
          pht_5_189 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_190 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15164) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_190 <= _pht_T_3;
        end else begin
          pht_5_190 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_191 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15167) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_191 <= _pht_T_3;
        end else begin
          pht_5_191 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_192 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15170) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_192 <= _pht_T_3;
        end else begin
          pht_5_192 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_193 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15173) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_193 <= _pht_T_3;
        end else begin
          pht_5_193 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_194 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15176) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_194 <= _pht_T_3;
        end else begin
          pht_5_194 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_195 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15179) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_195 <= _pht_T_3;
        end else begin
          pht_5_195 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_196 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15182) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_196 <= _pht_T_3;
        end else begin
          pht_5_196 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_197 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15185) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_197 <= _pht_T_3;
        end else begin
          pht_5_197 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_198 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15188) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_198 <= _pht_T_3;
        end else begin
          pht_5_198 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_199 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15191) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_199 <= _pht_T_3;
        end else begin
          pht_5_199 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_200 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15194) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_200 <= _pht_T_3;
        end else begin
          pht_5_200 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_201 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15197) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_201 <= _pht_T_3;
        end else begin
          pht_5_201 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_202 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15200) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_202 <= _pht_T_3;
        end else begin
          pht_5_202 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_203 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15203) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_203 <= _pht_T_3;
        end else begin
          pht_5_203 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_204 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15206) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_204 <= _pht_T_3;
        end else begin
          pht_5_204 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_205 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15209) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_205 <= _pht_T_3;
        end else begin
          pht_5_205 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_206 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15212) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_206 <= _pht_T_3;
        end else begin
          pht_5_206 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_207 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15215) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_207 <= _pht_T_3;
        end else begin
          pht_5_207 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_208 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15218) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_208 <= _pht_T_3;
        end else begin
          pht_5_208 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_209 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15221) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_209 <= _pht_T_3;
        end else begin
          pht_5_209 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_210 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15224) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_210 <= _pht_T_3;
        end else begin
          pht_5_210 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_211 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15227) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_211 <= _pht_T_3;
        end else begin
          pht_5_211 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_212 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15230) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_212 <= _pht_T_3;
        end else begin
          pht_5_212 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_213 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15233) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_213 <= _pht_T_3;
        end else begin
          pht_5_213 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_214 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15236) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_214 <= _pht_T_3;
        end else begin
          pht_5_214 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_215 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15239) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_215 <= _pht_T_3;
        end else begin
          pht_5_215 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_216 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15242) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_216 <= _pht_T_3;
        end else begin
          pht_5_216 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_217 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15245) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_217 <= _pht_T_3;
        end else begin
          pht_5_217 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_218 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15248) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_218 <= _pht_T_3;
        end else begin
          pht_5_218 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_219 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15251) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_219 <= _pht_T_3;
        end else begin
          pht_5_219 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_220 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15254) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_220 <= _pht_T_3;
        end else begin
          pht_5_220 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_221 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15257) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_221 <= _pht_T_3;
        end else begin
          pht_5_221 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_222 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15260) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_222 <= _pht_T_3;
        end else begin
          pht_5_222 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_223 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15263) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_223 <= _pht_T_3;
        end else begin
          pht_5_223 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_224 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15266) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_224 <= _pht_T_3;
        end else begin
          pht_5_224 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_225 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15269) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_225 <= _pht_T_3;
        end else begin
          pht_5_225 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_226 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15272) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_226 <= _pht_T_3;
        end else begin
          pht_5_226 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_227 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15275) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_227 <= _pht_T_3;
        end else begin
          pht_5_227 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_228 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15278) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_228 <= _pht_T_3;
        end else begin
          pht_5_228 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_229 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15281) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_229 <= _pht_T_3;
        end else begin
          pht_5_229 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_230 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15284) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_230 <= _pht_T_3;
        end else begin
          pht_5_230 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_231 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15287) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_231 <= _pht_T_3;
        end else begin
          pht_5_231 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_232 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15290) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_232 <= _pht_T_3;
        end else begin
          pht_5_232 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_233 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15293) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_233 <= _pht_T_3;
        end else begin
          pht_5_233 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_234 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15296) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_234 <= _pht_T_3;
        end else begin
          pht_5_234 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_235 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15299) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_235 <= _pht_T_3;
        end else begin
          pht_5_235 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_236 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15302) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_236 <= _pht_T_3;
        end else begin
          pht_5_236 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_237 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15305) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_237 <= _pht_T_3;
        end else begin
          pht_5_237 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_238 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15308) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_238 <= _pht_T_3;
        end else begin
          pht_5_238 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_239 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15311) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_239 <= _pht_T_3;
        end else begin
          pht_5_239 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_240 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15314) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_240 <= _pht_T_3;
        end else begin
          pht_5_240 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_241 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15317) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_241 <= _pht_T_3;
        end else begin
          pht_5_241 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_242 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15320) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_242 <= _pht_T_3;
        end else begin
          pht_5_242 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_243 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15323) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_243 <= _pht_T_3;
        end else begin
          pht_5_243 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_244 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15326) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_244 <= _pht_T_3;
        end else begin
          pht_5_244 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_245 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15329) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_245 <= _pht_T_3;
        end else begin
          pht_5_245 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_246 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15332) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_246 <= _pht_T_3;
        end else begin
          pht_5_246 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_247 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15335) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_247 <= _pht_T_3;
        end else begin
          pht_5_247 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_248 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15338) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_248 <= _pht_T_3;
        end else begin
          pht_5_248 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_249 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15341) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_249 <= _pht_T_3;
        end else begin
          pht_5_249 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_250 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15344) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_250 <= _pht_T_3;
        end else begin
          pht_5_250 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_251 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15347) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_251 <= _pht_T_3;
        end else begin
          pht_5_251 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_252 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15350) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_252 <= _pht_T_3;
        end else begin
          pht_5_252 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_253 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15353) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_253 <= _pht_T_3;
        end else begin
          pht_5_253 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_254 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15356) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_254 <= _pht_T_3;
        end else begin
          pht_5_254 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_5_255 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18176 & _GEN_15359) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_5_255 <= _pht_T_3;
        end else begin
          pht_5_255 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_0 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15361) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_0 <= _pht_T_3;
        end else begin
          pht_6_0 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_1 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14659) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_1 <= _pht_T_3;
        end else begin
          pht_6_1 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_2 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14661) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_2 <= _pht_T_3;
        end else begin
          pht_6_2 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_3 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14663) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_3 <= _pht_T_3;
        end else begin
          pht_6_3 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_4 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14665) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_4 <= _pht_T_3;
        end else begin
          pht_6_4 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_5 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14667) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_5 <= _pht_T_3;
        end else begin
          pht_6_5 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_6 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14669) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_6 <= _pht_T_3;
        end else begin
          pht_6_6 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_7 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14671) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_7 <= _pht_T_3;
        end else begin
          pht_6_7 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_8 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14673) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_8 <= _pht_T_3;
        end else begin
          pht_6_8 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_9 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14675) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_9 <= _pht_T_3;
        end else begin
          pht_6_9 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_10 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14677) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_10 <= _pht_T_3;
        end else begin
          pht_6_10 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_11 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14679) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_11 <= _pht_T_3;
        end else begin
          pht_6_11 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_12 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14681) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_12 <= _pht_T_3;
        end else begin
          pht_6_12 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_13 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14683) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_13 <= _pht_T_3;
        end else begin
          pht_6_13 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_14 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14685) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_14 <= _pht_T_3;
        end else begin
          pht_6_14 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_15 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14687) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_15 <= _pht_T_3;
        end else begin
          pht_6_15 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_16 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14689) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_16 <= _pht_T_3;
        end else begin
          pht_6_16 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_17 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14691) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_17 <= _pht_T_3;
        end else begin
          pht_6_17 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_18 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14693) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_18 <= _pht_T_3;
        end else begin
          pht_6_18 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_19 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14695) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_19 <= _pht_T_3;
        end else begin
          pht_6_19 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_20 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14697) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_20 <= _pht_T_3;
        end else begin
          pht_6_20 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_21 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14699) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_21 <= _pht_T_3;
        end else begin
          pht_6_21 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_22 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14701) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_22 <= _pht_T_3;
        end else begin
          pht_6_22 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_23 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14703) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_23 <= _pht_T_3;
        end else begin
          pht_6_23 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_24 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14705) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_24 <= _pht_T_3;
        end else begin
          pht_6_24 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_25 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14707) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_25 <= _pht_T_3;
        end else begin
          pht_6_25 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_26 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14709) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_26 <= _pht_T_3;
        end else begin
          pht_6_26 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_27 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14711) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_27 <= _pht_T_3;
        end else begin
          pht_6_27 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_28 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14713) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_28 <= _pht_T_3;
        end else begin
          pht_6_28 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_29 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14715) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_29 <= _pht_T_3;
        end else begin
          pht_6_29 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_30 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14717) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_30 <= _pht_T_3;
        end else begin
          pht_6_30 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_31 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14719) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_31 <= _pht_T_3;
        end else begin
          pht_6_31 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_32 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14721) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_32 <= _pht_T_3;
        end else begin
          pht_6_32 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_33 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14723) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_33 <= _pht_T_3;
        end else begin
          pht_6_33 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_34 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14725) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_34 <= _pht_T_3;
        end else begin
          pht_6_34 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_35 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14727) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_35 <= _pht_T_3;
        end else begin
          pht_6_35 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_36 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14729) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_36 <= _pht_T_3;
        end else begin
          pht_6_36 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_37 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14731) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_37 <= _pht_T_3;
        end else begin
          pht_6_37 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_38 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14733) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_38 <= _pht_T_3;
        end else begin
          pht_6_38 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_39 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14735) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_39 <= _pht_T_3;
        end else begin
          pht_6_39 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_40 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14737) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_40 <= _pht_T_3;
        end else begin
          pht_6_40 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_41 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14739) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_41 <= _pht_T_3;
        end else begin
          pht_6_41 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_42 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14741) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_42 <= _pht_T_3;
        end else begin
          pht_6_42 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_43 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14743) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_43 <= _pht_T_3;
        end else begin
          pht_6_43 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_44 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14745) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_44 <= _pht_T_3;
        end else begin
          pht_6_44 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_45 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14747) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_45 <= _pht_T_3;
        end else begin
          pht_6_45 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_46 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14749) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_46 <= _pht_T_3;
        end else begin
          pht_6_46 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_47 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14751) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_47 <= _pht_T_3;
        end else begin
          pht_6_47 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_48 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14753) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_48 <= _pht_T_3;
        end else begin
          pht_6_48 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_49 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14755) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_49 <= _pht_T_3;
        end else begin
          pht_6_49 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_50 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14757) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_50 <= _pht_T_3;
        end else begin
          pht_6_50 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_51 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14759) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_51 <= _pht_T_3;
        end else begin
          pht_6_51 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_52 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14761) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_52 <= _pht_T_3;
        end else begin
          pht_6_52 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_53 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14763) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_53 <= _pht_T_3;
        end else begin
          pht_6_53 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_54 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14765) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_54 <= _pht_T_3;
        end else begin
          pht_6_54 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_55 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14767) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_55 <= _pht_T_3;
        end else begin
          pht_6_55 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_56 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14769) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_56 <= _pht_T_3;
        end else begin
          pht_6_56 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_57 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14771) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_57 <= _pht_T_3;
        end else begin
          pht_6_57 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_58 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14773) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_58 <= _pht_T_3;
        end else begin
          pht_6_58 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_59 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14775) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_59 <= _pht_T_3;
        end else begin
          pht_6_59 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_60 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14777) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_60 <= _pht_T_3;
        end else begin
          pht_6_60 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_61 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14779) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_61 <= _pht_T_3;
        end else begin
          pht_6_61 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_62 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14781) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_62 <= _pht_T_3;
        end else begin
          pht_6_62 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_63 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14783) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_63 <= _pht_T_3;
        end else begin
          pht_6_63 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_64 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14786) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_64 <= _pht_T_3;
        end else begin
          pht_6_64 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_65 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14789) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_65 <= _pht_T_3;
        end else begin
          pht_6_65 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_66 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14792) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_66 <= _pht_T_3;
        end else begin
          pht_6_66 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_67 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14795) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_67 <= _pht_T_3;
        end else begin
          pht_6_67 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_68 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14798) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_68 <= _pht_T_3;
        end else begin
          pht_6_68 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_69 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14801) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_69 <= _pht_T_3;
        end else begin
          pht_6_69 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_70 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14804) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_70 <= _pht_T_3;
        end else begin
          pht_6_70 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_71 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14807) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_71 <= _pht_T_3;
        end else begin
          pht_6_71 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_72 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14810) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_72 <= _pht_T_3;
        end else begin
          pht_6_72 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_73 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14813) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_73 <= _pht_T_3;
        end else begin
          pht_6_73 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_74 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14816) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_74 <= _pht_T_3;
        end else begin
          pht_6_74 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_75 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14819) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_75 <= _pht_T_3;
        end else begin
          pht_6_75 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_76 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14822) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_76 <= _pht_T_3;
        end else begin
          pht_6_76 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_77 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14825) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_77 <= _pht_T_3;
        end else begin
          pht_6_77 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_78 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14828) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_78 <= _pht_T_3;
        end else begin
          pht_6_78 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_79 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14831) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_79 <= _pht_T_3;
        end else begin
          pht_6_79 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_80 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14834) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_80 <= _pht_T_3;
        end else begin
          pht_6_80 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_81 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14837) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_81 <= _pht_T_3;
        end else begin
          pht_6_81 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_82 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14840) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_82 <= _pht_T_3;
        end else begin
          pht_6_82 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_83 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14843) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_83 <= _pht_T_3;
        end else begin
          pht_6_83 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_84 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14846) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_84 <= _pht_T_3;
        end else begin
          pht_6_84 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_85 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14849) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_85 <= _pht_T_3;
        end else begin
          pht_6_85 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_86 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14852) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_86 <= _pht_T_3;
        end else begin
          pht_6_86 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_87 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14855) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_87 <= _pht_T_3;
        end else begin
          pht_6_87 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_88 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14858) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_88 <= _pht_T_3;
        end else begin
          pht_6_88 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_89 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14861) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_89 <= _pht_T_3;
        end else begin
          pht_6_89 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_90 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14864) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_90 <= _pht_T_3;
        end else begin
          pht_6_90 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_91 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14867) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_91 <= _pht_T_3;
        end else begin
          pht_6_91 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_92 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14870) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_92 <= _pht_T_3;
        end else begin
          pht_6_92 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_93 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14873) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_93 <= _pht_T_3;
        end else begin
          pht_6_93 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_94 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14876) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_94 <= _pht_T_3;
        end else begin
          pht_6_94 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_95 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14879) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_95 <= _pht_T_3;
        end else begin
          pht_6_95 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_96 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14882) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_96 <= _pht_T_3;
        end else begin
          pht_6_96 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_97 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14885) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_97 <= _pht_T_3;
        end else begin
          pht_6_97 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_98 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14888) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_98 <= _pht_T_3;
        end else begin
          pht_6_98 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_99 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14891) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_99 <= _pht_T_3;
        end else begin
          pht_6_99 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_100 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14894) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_100 <= _pht_T_3;
        end else begin
          pht_6_100 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_101 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14897) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_101 <= _pht_T_3;
        end else begin
          pht_6_101 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_102 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14900) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_102 <= _pht_T_3;
        end else begin
          pht_6_102 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_103 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14903) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_103 <= _pht_T_3;
        end else begin
          pht_6_103 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_104 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14906) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_104 <= _pht_T_3;
        end else begin
          pht_6_104 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_105 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14909) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_105 <= _pht_T_3;
        end else begin
          pht_6_105 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_106 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14912) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_106 <= _pht_T_3;
        end else begin
          pht_6_106 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_107 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14915) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_107 <= _pht_T_3;
        end else begin
          pht_6_107 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_108 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14918) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_108 <= _pht_T_3;
        end else begin
          pht_6_108 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_109 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14921) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_109 <= _pht_T_3;
        end else begin
          pht_6_109 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_110 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14924) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_110 <= _pht_T_3;
        end else begin
          pht_6_110 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_111 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14927) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_111 <= _pht_T_3;
        end else begin
          pht_6_111 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_112 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14930) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_112 <= _pht_T_3;
        end else begin
          pht_6_112 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_113 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14933) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_113 <= _pht_T_3;
        end else begin
          pht_6_113 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_114 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14936) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_114 <= _pht_T_3;
        end else begin
          pht_6_114 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_115 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14939) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_115 <= _pht_T_3;
        end else begin
          pht_6_115 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_116 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14942) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_116 <= _pht_T_3;
        end else begin
          pht_6_116 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_117 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14945) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_117 <= _pht_T_3;
        end else begin
          pht_6_117 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_118 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14948) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_118 <= _pht_T_3;
        end else begin
          pht_6_118 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_119 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14951) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_119 <= _pht_T_3;
        end else begin
          pht_6_119 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_120 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14954) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_120 <= _pht_T_3;
        end else begin
          pht_6_120 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_121 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14957) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_121 <= _pht_T_3;
        end else begin
          pht_6_121 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_122 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14960) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_122 <= _pht_T_3;
        end else begin
          pht_6_122 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_123 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14963) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_123 <= _pht_T_3;
        end else begin
          pht_6_123 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_124 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14966) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_124 <= _pht_T_3;
        end else begin
          pht_6_124 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_125 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14969) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_125 <= _pht_T_3;
        end else begin
          pht_6_125 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_126 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14972) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_126 <= _pht_T_3;
        end else begin
          pht_6_126 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_127 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14975) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_127 <= _pht_T_3;
        end else begin
          pht_6_127 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_128 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14978) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_128 <= _pht_T_3;
        end else begin
          pht_6_128 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_129 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14981) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_129 <= _pht_T_3;
        end else begin
          pht_6_129 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_130 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14984) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_130 <= _pht_T_3;
        end else begin
          pht_6_130 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_131 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14987) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_131 <= _pht_T_3;
        end else begin
          pht_6_131 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_132 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14990) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_132 <= _pht_T_3;
        end else begin
          pht_6_132 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_133 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14993) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_133 <= _pht_T_3;
        end else begin
          pht_6_133 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_134 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14996) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_134 <= _pht_T_3;
        end else begin
          pht_6_134 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_135 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_14999) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_135 <= _pht_T_3;
        end else begin
          pht_6_135 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_136 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15002) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_136 <= _pht_T_3;
        end else begin
          pht_6_136 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_137 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15005) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_137 <= _pht_T_3;
        end else begin
          pht_6_137 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_138 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15008) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_138 <= _pht_T_3;
        end else begin
          pht_6_138 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_139 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15011) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_139 <= _pht_T_3;
        end else begin
          pht_6_139 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_140 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15014) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_140 <= _pht_T_3;
        end else begin
          pht_6_140 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_141 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15017) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_141 <= _pht_T_3;
        end else begin
          pht_6_141 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_142 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15020) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_142 <= _pht_T_3;
        end else begin
          pht_6_142 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_143 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15023) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_143 <= _pht_T_3;
        end else begin
          pht_6_143 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_144 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15026) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_144 <= _pht_T_3;
        end else begin
          pht_6_144 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_145 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15029) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_145 <= _pht_T_3;
        end else begin
          pht_6_145 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_146 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15032) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_146 <= _pht_T_3;
        end else begin
          pht_6_146 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_147 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15035) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_147 <= _pht_T_3;
        end else begin
          pht_6_147 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_148 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15038) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_148 <= _pht_T_3;
        end else begin
          pht_6_148 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_149 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15041) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_149 <= _pht_T_3;
        end else begin
          pht_6_149 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_150 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15044) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_150 <= _pht_T_3;
        end else begin
          pht_6_150 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_151 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15047) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_151 <= _pht_T_3;
        end else begin
          pht_6_151 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_152 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15050) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_152 <= _pht_T_3;
        end else begin
          pht_6_152 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_153 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15053) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_153 <= _pht_T_3;
        end else begin
          pht_6_153 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_154 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15056) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_154 <= _pht_T_3;
        end else begin
          pht_6_154 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_155 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15059) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_155 <= _pht_T_3;
        end else begin
          pht_6_155 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_156 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15062) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_156 <= _pht_T_3;
        end else begin
          pht_6_156 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_157 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15065) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_157 <= _pht_T_3;
        end else begin
          pht_6_157 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_158 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15068) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_158 <= _pht_T_3;
        end else begin
          pht_6_158 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_159 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15071) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_159 <= _pht_T_3;
        end else begin
          pht_6_159 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_160 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15074) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_160 <= _pht_T_3;
        end else begin
          pht_6_160 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_161 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15077) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_161 <= _pht_T_3;
        end else begin
          pht_6_161 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_162 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15080) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_162 <= _pht_T_3;
        end else begin
          pht_6_162 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_163 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15083) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_163 <= _pht_T_3;
        end else begin
          pht_6_163 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_164 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15086) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_164 <= _pht_T_3;
        end else begin
          pht_6_164 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_165 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15089) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_165 <= _pht_T_3;
        end else begin
          pht_6_165 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_166 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15092) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_166 <= _pht_T_3;
        end else begin
          pht_6_166 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_167 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15095) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_167 <= _pht_T_3;
        end else begin
          pht_6_167 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_168 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15098) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_168 <= _pht_T_3;
        end else begin
          pht_6_168 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_169 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15101) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_169 <= _pht_T_3;
        end else begin
          pht_6_169 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_170 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15104) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_170 <= _pht_T_3;
        end else begin
          pht_6_170 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_171 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15107) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_171 <= _pht_T_3;
        end else begin
          pht_6_171 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_172 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15110) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_172 <= _pht_T_3;
        end else begin
          pht_6_172 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_173 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15113) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_173 <= _pht_T_3;
        end else begin
          pht_6_173 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_174 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15116) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_174 <= _pht_T_3;
        end else begin
          pht_6_174 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_175 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15119) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_175 <= _pht_T_3;
        end else begin
          pht_6_175 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_176 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15122) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_176 <= _pht_T_3;
        end else begin
          pht_6_176 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_177 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15125) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_177 <= _pht_T_3;
        end else begin
          pht_6_177 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_178 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15128) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_178 <= _pht_T_3;
        end else begin
          pht_6_178 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_179 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15131) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_179 <= _pht_T_3;
        end else begin
          pht_6_179 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_180 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15134) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_180 <= _pht_T_3;
        end else begin
          pht_6_180 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_181 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15137) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_181 <= _pht_T_3;
        end else begin
          pht_6_181 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_182 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15140) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_182 <= _pht_T_3;
        end else begin
          pht_6_182 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_183 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15143) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_183 <= _pht_T_3;
        end else begin
          pht_6_183 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_184 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15146) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_184 <= _pht_T_3;
        end else begin
          pht_6_184 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_185 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15149) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_185 <= _pht_T_3;
        end else begin
          pht_6_185 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_186 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15152) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_186 <= _pht_T_3;
        end else begin
          pht_6_186 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_187 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15155) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_187 <= _pht_T_3;
        end else begin
          pht_6_187 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_188 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15158) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_188 <= _pht_T_3;
        end else begin
          pht_6_188 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_189 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15161) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_189 <= _pht_T_3;
        end else begin
          pht_6_189 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_190 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15164) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_190 <= _pht_T_3;
        end else begin
          pht_6_190 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_191 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15167) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_191 <= _pht_T_3;
        end else begin
          pht_6_191 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_192 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15170) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_192 <= _pht_T_3;
        end else begin
          pht_6_192 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_193 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15173) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_193 <= _pht_T_3;
        end else begin
          pht_6_193 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_194 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15176) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_194 <= _pht_T_3;
        end else begin
          pht_6_194 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_195 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15179) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_195 <= _pht_T_3;
        end else begin
          pht_6_195 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_196 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15182) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_196 <= _pht_T_3;
        end else begin
          pht_6_196 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_197 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15185) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_197 <= _pht_T_3;
        end else begin
          pht_6_197 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_198 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15188) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_198 <= _pht_T_3;
        end else begin
          pht_6_198 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_199 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15191) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_199 <= _pht_T_3;
        end else begin
          pht_6_199 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_200 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15194) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_200 <= _pht_T_3;
        end else begin
          pht_6_200 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_201 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15197) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_201 <= _pht_T_3;
        end else begin
          pht_6_201 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_202 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15200) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_202 <= _pht_T_3;
        end else begin
          pht_6_202 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_203 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15203) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_203 <= _pht_T_3;
        end else begin
          pht_6_203 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_204 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15206) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_204 <= _pht_T_3;
        end else begin
          pht_6_204 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_205 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15209) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_205 <= _pht_T_3;
        end else begin
          pht_6_205 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_206 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15212) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_206 <= _pht_T_3;
        end else begin
          pht_6_206 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_207 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15215) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_207 <= _pht_T_3;
        end else begin
          pht_6_207 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_208 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15218) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_208 <= _pht_T_3;
        end else begin
          pht_6_208 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_209 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15221) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_209 <= _pht_T_3;
        end else begin
          pht_6_209 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_210 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15224) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_210 <= _pht_T_3;
        end else begin
          pht_6_210 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_211 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15227) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_211 <= _pht_T_3;
        end else begin
          pht_6_211 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_212 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15230) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_212 <= _pht_T_3;
        end else begin
          pht_6_212 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_213 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15233) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_213 <= _pht_T_3;
        end else begin
          pht_6_213 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_214 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15236) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_214 <= _pht_T_3;
        end else begin
          pht_6_214 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_215 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15239) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_215 <= _pht_T_3;
        end else begin
          pht_6_215 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_216 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15242) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_216 <= _pht_T_3;
        end else begin
          pht_6_216 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_217 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15245) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_217 <= _pht_T_3;
        end else begin
          pht_6_217 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_218 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15248) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_218 <= _pht_T_3;
        end else begin
          pht_6_218 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_219 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15251) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_219 <= _pht_T_3;
        end else begin
          pht_6_219 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_220 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15254) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_220 <= _pht_T_3;
        end else begin
          pht_6_220 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_221 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15257) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_221 <= _pht_T_3;
        end else begin
          pht_6_221 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_222 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15260) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_222 <= _pht_T_3;
        end else begin
          pht_6_222 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_223 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15263) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_223 <= _pht_T_3;
        end else begin
          pht_6_223 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_224 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15266) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_224 <= _pht_T_3;
        end else begin
          pht_6_224 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_225 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15269) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_225 <= _pht_T_3;
        end else begin
          pht_6_225 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_226 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15272) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_226 <= _pht_T_3;
        end else begin
          pht_6_226 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_227 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15275) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_227 <= _pht_T_3;
        end else begin
          pht_6_227 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_228 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15278) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_228 <= _pht_T_3;
        end else begin
          pht_6_228 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_229 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15281) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_229 <= _pht_T_3;
        end else begin
          pht_6_229 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_230 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15284) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_230 <= _pht_T_3;
        end else begin
          pht_6_230 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_231 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15287) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_231 <= _pht_T_3;
        end else begin
          pht_6_231 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_232 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15290) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_232 <= _pht_T_3;
        end else begin
          pht_6_232 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_233 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15293) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_233 <= _pht_T_3;
        end else begin
          pht_6_233 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_234 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15296) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_234 <= _pht_T_3;
        end else begin
          pht_6_234 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_235 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15299) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_235 <= _pht_T_3;
        end else begin
          pht_6_235 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_236 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15302) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_236 <= _pht_T_3;
        end else begin
          pht_6_236 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_237 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15305) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_237 <= _pht_T_3;
        end else begin
          pht_6_237 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_238 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15308) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_238 <= _pht_T_3;
        end else begin
          pht_6_238 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_239 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15311) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_239 <= _pht_T_3;
        end else begin
          pht_6_239 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_240 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15314) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_240 <= _pht_T_3;
        end else begin
          pht_6_240 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_241 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15317) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_241 <= _pht_T_3;
        end else begin
          pht_6_241 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_242 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15320) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_242 <= _pht_T_3;
        end else begin
          pht_6_242 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_243 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15323) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_243 <= _pht_T_3;
        end else begin
          pht_6_243 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_244 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15326) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_244 <= _pht_T_3;
        end else begin
          pht_6_244 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_245 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15329) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_245 <= _pht_T_3;
        end else begin
          pht_6_245 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_246 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15332) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_246 <= _pht_T_3;
        end else begin
          pht_6_246 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_247 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15335) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_247 <= _pht_T_3;
        end else begin
          pht_6_247 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_248 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15338) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_248 <= _pht_T_3;
        end else begin
          pht_6_248 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_249 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15341) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_249 <= _pht_T_3;
        end else begin
          pht_6_249 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_250 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15344) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_250 <= _pht_T_3;
        end else begin
          pht_6_250 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_251 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15347) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_251 <= _pht_T_3;
        end else begin
          pht_6_251 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_252 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15350) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_252 <= _pht_T_3;
        end else begin
          pht_6_252 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_253 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15353) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_253 <= _pht_T_3;
        end else begin
          pht_6_253 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_254 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15356) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_254 <= _pht_T_3;
        end else begin
          pht_6_254 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_6_255 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_18880 & _GEN_15359) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_6_255 <= _pht_T_3;
        end else begin
          pht_6_255 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_0 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15361) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_0 <= _pht_T_3;
        end else begin
          pht_7_0 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_1 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14659) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_1 <= _pht_T_3;
        end else begin
          pht_7_1 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_2 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14661) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_2 <= _pht_T_3;
        end else begin
          pht_7_2 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_3 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14663) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_3 <= _pht_T_3;
        end else begin
          pht_7_3 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_4 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14665) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_4 <= _pht_T_3;
        end else begin
          pht_7_4 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_5 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14667) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_5 <= _pht_T_3;
        end else begin
          pht_7_5 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_6 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14669) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_6 <= _pht_T_3;
        end else begin
          pht_7_6 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_7 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14671) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_7 <= _pht_T_3;
        end else begin
          pht_7_7 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_8 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14673) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_8 <= _pht_T_3;
        end else begin
          pht_7_8 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_9 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14675) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_9 <= _pht_T_3;
        end else begin
          pht_7_9 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_10 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14677) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_10 <= _pht_T_3;
        end else begin
          pht_7_10 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_11 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14679) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_11 <= _pht_T_3;
        end else begin
          pht_7_11 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_12 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14681) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_12 <= _pht_T_3;
        end else begin
          pht_7_12 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_13 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14683) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_13 <= _pht_T_3;
        end else begin
          pht_7_13 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_14 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14685) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_14 <= _pht_T_3;
        end else begin
          pht_7_14 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_15 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14687) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_15 <= _pht_T_3;
        end else begin
          pht_7_15 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_16 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14689) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_16 <= _pht_T_3;
        end else begin
          pht_7_16 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_17 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14691) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_17 <= _pht_T_3;
        end else begin
          pht_7_17 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_18 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14693) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_18 <= _pht_T_3;
        end else begin
          pht_7_18 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_19 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14695) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_19 <= _pht_T_3;
        end else begin
          pht_7_19 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_20 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14697) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_20 <= _pht_T_3;
        end else begin
          pht_7_20 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_21 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14699) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_21 <= _pht_T_3;
        end else begin
          pht_7_21 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_22 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14701) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_22 <= _pht_T_3;
        end else begin
          pht_7_22 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_23 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14703) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_23 <= _pht_T_3;
        end else begin
          pht_7_23 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_24 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14705) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_24 <= _pht_T_3;
        end else begin
          pht_7_24 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_25 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14707) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_25 <= _pht_T_3;
        end else begin
          pht_7_25 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_26 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14709) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_26 <= _pht_T_3;
        end else begin
          pht_7_26 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_27 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14711) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_27 <= _pht_T_3;
        end else begin
          pht_7_27 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_28 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14713) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_28 <= _pht_T_3;
        end else begin
          pht_7_28 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_29 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14715) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_29 <= _pht_T_3;
        end else begin
          pht_7_29 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_30 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14717) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_30 <= _pht_T_3;
        end else begin
          pht_7_30 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_31 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14719) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_31 <= _pht_T_3;
        end else begin
          pht_7_31 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_32 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14721) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_32 <= _pht_T_3;
        end else begin
          pht_7_32 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_33 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14723) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_33 <= _pht_T_3;
        end else begin
          pht_7_33 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_34 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14725) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_34 <= _pht_T_3;
        end else begin
          pht_7_34 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_35 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14727) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_35 <= _pht_T_3;
        end else begin
          pht_7_35 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_36 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14729) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_36 <= _pht_T_3;
        end else begin
          pht_7_36 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_37 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14731) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_37 <= _pht_T_3;
        end else begin
          pht_7_37 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_38 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14733) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_38 <= _pht_T_3;
        end else begin
          pht_7_38 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_39 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14735) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_39 <= _pht_T_3;
        end else begin
          pht_7_39 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_40 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14737) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_40 <= _pht_T_3;
        end else begin
          pht_7_40 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_41 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14739) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_41 <= _pht_T_3;
        end else begin
          pht_7_41 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_42 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14741) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_42 <= _pht_T_3;
        end else begin
          pht_7_42 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_43 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14743) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_43 <= _pht_T_3;
        end else begin
          pht_7_43 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_44 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14745) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_44 <= _pht_T_3;
        end else begin
          pht_7_44 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_45 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14747) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_45 <= _pht_T_3;
        end else begin
          pht_7_45 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_46 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14749) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_46 <= _pht_T_3;
        end else begin
          pht_7_46 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_47 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14751) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_47 <= _pht_T_3;
        end else begin
          pht_7_47 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_48 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14753) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_48 <= _pht_T_3;
        end else begin
          pht_7_48 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_49 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14755) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_49 <= _pht_T_3;
        end else begin
          pht_7_49 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_50 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14757) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_50 <= _pht_T_3;
        end else begin
          pht_7_50 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_51 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14759) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_51 <= _pht_T_3;
        end else begin
          pht_7_51 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_52 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14761) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_52 <= _pht_T_3;
        end else begin
          pht_7_52 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_53 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14763) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_53 <= _pht_T_3;
        end else begin
          pht_7_53 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_54 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14765) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_54 <= _pht_T_3;
        end else begin
          pht_7_54 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_55 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14767) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_55 <= _pht_T_3;
        end else begin
          pht_7_55 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_56 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14769) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_56 <= _pht_T_3;
        end else begin
          pht_7_56 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_57 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14771) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_57 <= _pht_T_3;
        end else begin
          pht_7_57 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_58 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14773) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_58 <= _pht_T_3;
        end else begin
          pht_7_58 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_59 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14775) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_59 <= _pht_T_3;
        end else begin
          pht_7_59 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_60 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14777) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_60 <= _pht_T_3;
        end else begin
          pht_7_60 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_61 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14779) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_61 <= _pht_T_3;
        end else begin
          pht_7_61 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_62 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14781) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_62 <= _pht_T_3;
        end else begin
          pht_7_62 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_63 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14783) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_63 <= _pht_T_3;
        end else begin
          pht_7_63 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_64 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14786) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_64 <= _pht_T_3;
        end else begin
          pht_7_64 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_65 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14789) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_65 <= _pht_T_3;
        end else begin
          pht_7_65 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_66 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14792) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_66 <= _pht_T_3;
        end else begin
          pht_7_66 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_67 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14795) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_67 <= _pht_T_3;
        end else begin
          pht_7_67 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_68 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14798) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_68 <= _pht_T_3;
        end else begin
          pht_7_68 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_69 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14801) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_69 <= _pht_T_3;
        end else begin
          pht_7_69 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_70 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14804) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_70 <= _pht_T_3;
        end else begin
          pht_7_70 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_71 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14807) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_71 <= _pht_T_3;
        end else begin
          pht_7_71 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_72 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14810) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_72 <= _pht_T_3;
        end else begin
          pht_7_72 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_73 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14813) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_73 <= _pht_T_3;
        end else begin
          pht_7_73 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_74 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14816) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_74 <= _pht_T_3;
        end else begin
          pht_7_74 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_75 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14819) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_75 <= _pht_T_3;
        end else begin
          pht_7_75 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_76 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14822) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_76 <= _pht_T_3;
        end else begin
          pht_7_76 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_77 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14825) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_77 <= _pht_T_3;
        end else begin
          pht_7_77 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_78 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14828) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_78 <= _pht_T_3;
        end else begin
          pht_7_78 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_79 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14831) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_79 <= _pht_T_3;
        end else begin
          pht_7_79 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_80 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14834) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_80 <= _pht_T_3;
        end else begin
          pht_7_80 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_81 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14837) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_81 <= _pht_T_3;
        end else begin
          pht_7_81 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_82 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14840) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_82 <= _pht_T_3;
        end else begin
          pht_7_82 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_83 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14843) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_83 <= _pht_T_3;
        end else begin
          pht_7_83 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_84 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14846) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_84 <= _pht_T_3;
        end else begin
          pht_7_84 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_85 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14849) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_85 <= _pht_T_3;
        end else begin
          pht_7_85 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_86 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14852) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_86 <= _pht_T_3;
        end else begin
          pht_7_86 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_87 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14855) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_87 <= _pht_T_3;
        end else begin
          pht_7_87 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_88 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14858) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_88 <= _pht_T_3;
        end else begin
          pht_7_88 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_89 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14861) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_89 <= _pht_T_3;
        end else begin
          pht_7_89 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_90 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14864) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_90 <= _pht_T_3;
        end else begin
          pht_7_90 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_91 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14867) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_91 <= _pht_T_3;
        end else begin
          pht_7_91 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_92 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14870) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_92 <= _pht_T_3;
        end else begin
          pht_7_92 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_93 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14873) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_93 <= _pht_T_3;
        end else begin
          pht_7_93 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_94 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14876) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_94 <= _pht_T_3;
        end else begin
          pht_7_94 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_95 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14879) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_95 <= _pht_T_3;
        end else begin
          pht_7_95 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_96 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14882) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_96 <= _pht_T_3;
        end else begin
          pht_7_96 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_97 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14885) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_97 <= _pht_T_3;
        end else begin
          pht_7_97 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_98 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14888) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_98 <= _pht_T_3;
        end else begin
          pht_7_98 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_99 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14891) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_99 <= _pht_T_3;
        end else begin
          pht_7_99 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_100 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14894) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_100 <= _pht_T_3;
        end else begin
          pht_7_100 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_101 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14897) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_101 <= _pht_T_3;
        end else begin
          pht_7_101 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_102 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14900) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_102 <= _pht_T_3;
        end else begin
          pht_7_102 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_103 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14903) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_103 <= _pht_T_3;
        end else begin
          pht_7_103 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_104 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14906) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_104 <= _pht_T_3;
        end else begin
          pht_7_104 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_105 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14909) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_105 <= _pht_T_3;
        end else begin
          pht_7_105 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_106 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14912) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_106 <= _pht_T_3;
        end else begin
          pht_7_106 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_107 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14915) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_107 <= _pht_T_3;
        end else begin
          pht_7_107 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_108 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14918) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_108 <= _pht_T_3;
        end else begin
          pht_7_108 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_109 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14921) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_109 <= _pht_T_3;
        end else begin
          pht_7_109 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_110 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14924) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_110 <= _pht_T_3;
        end else begin
          pht_7_110 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_111 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14927) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_111 <= _pht_T_3;
        end else begin
          pht_7_111 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_112 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14930) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_112 <= _pht_T_3;
        end else begin
          pht_7_112 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_113 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14933) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_113 <= _pht_T_3;
        end else begin
          pht_7_113 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_114 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14936) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_114 <= _pht_T_3;
        end else begin
          pht_7_114 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_115 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14939) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_115 <= _pht_T_3;
        end else begin
          pht_7_115 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_116 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14942) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_116 <= _pht_T_3;
        end else begin
          pht_7_116 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_117 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14945) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_117 <= _pht_T_3;
        end else begin
          pht_7_117 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_118 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14948) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_118 <= _pht_T_3;
        end else begin
          pht_7_118 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_119 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14951) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_119 <= _pht_T_3;
        end else begin
          pht_7_119 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_120 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14954) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_120 <= _pht_T_3;
        end else begin
          pht_7_120 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_121 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14957) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_121 <= _pht_T_3;
        end else begin
          pht_7_121 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_122 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14960) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_122 <= _pht_T_3;
        end else begin
          pht_7_122 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_123 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14963) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_123 <= _pht_T_3;
        end else begin
          pht_7_123 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_124 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14966) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_124 <= _pht_T_3;
        end else begin
          pht_7_124 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_125 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14969) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_125 <= _pht_T_3;
        end else begin
          pht_7_125 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_126 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14972) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_126 <= _pht_T_3;
        end else begin
          pht_7_126 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_127 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14975) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_127 <= _pht_T_3;
        end else begin
          pht_7_127 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_128 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14978) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_128 <= _pht_T_3;
        end else begin
          pht_7_128 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_129 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14981) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_129 <= _pht_T_3;
        end else begin
          pht_7_129 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_130 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14984) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_130 <= _pht_T_3;
        end else begin
          pht_7_130 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_131 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14987) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_131 <= _pht_T_3;
        end else begin
          pht_7_131 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_132 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14990) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_132 <= _pht_T_3;
        end else begin
          pht_7_132 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_133 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14993) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_133 <= _pht_T_3;
        end else begin
          pht_7_133 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_134 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14996) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_134 <= _pht_T_3;
        end else begin
          pht_7_134 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_135 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_14999) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_135 <= _pht_T_3;
        end else begin
          pht_7_135 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_136 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15002) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_136 <= _pht_T_3;
        end else begin
          pht_7_136 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_137 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15005) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_137 <= _pht_T_3;
        end else begin
          pht_7_137 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_138 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15008) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_138 <= _pht_T_3;
        end else begin
          pht_7_138 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_139 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15011) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_139 <= _pht_T_3;
        end else begin
          pht_7_139 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_140 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15014) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_140 <= _pht_T_3;
        end else begin
          pht_7_140 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_141 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15017) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_141 <= _pht_T_3;
        end else begin
          pht_7_141 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_142 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15020) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_142 <= _pht_T_3;
        end else begin
          pht_7_142 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_143 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15023) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_143 <= _pht_T_3;
        end else begin
          pht_7_143 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_144 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15026) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_144 <= _pht_T_3;
        end else begin
          pht_7_144 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_145 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15029) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_145 <= _pht_T_3;
        end else begin
          pht_7_145 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_146 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15032) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_146 <= _pht_T_3;
        end else begin
          pht_7_146 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_147 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15035) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_147 <= _pht_T_3;
        end else begin
          pht_7_147 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_148 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15038) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_148 <= _pht_T_3;
        end else begin
          pht_7_148 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_149 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15041) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_149 <= _pht_T_3;
        end else begin
          pht_7_149 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_150 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15044) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_150 <= _pht_T_3;
        end else begin
          pht_7_150 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_151 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15047) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_151 <= _pht_T_3;
        end else begin
          pht_7_151 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_152 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15050) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_152 <= _pht_T_3;
        end else begin
          pht_7_152 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_153 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15053) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_153 <= _pht_T_3;
        end else begin
          pht_7_153 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_154 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15056) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_154 <= _pht_T_3;
        end else begin
          pht_7_154 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_155 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15059) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_155 <= _pht_T_3;
        end else begin
          pht_7_155 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_156 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15062) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_156 <= _pht_T_3;
        end else begin
          pht_7_156 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_157 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15065) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_157 <= _pht_T_3;
        end else begin
          pht_7_157 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_158 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15068) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_158 <= _pht_T_3;
        end else begin
          pht_7_158 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_159 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15071) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_159 <= _pht_T_3;
        end else begin
          pht_7_159 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_160 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15074) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_160 <= _pht_T_3;
        end else begin
          pht_7_160 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_161 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15077) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_161 <= _pht_T_3;
        end else begin
          pht_7_161 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_162 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15080) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_162 <= _pht_T_3;
        end else begin
          pht_7_162 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_163 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15083) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_163 <= _pht_T_3;
        end else begin
          pht_7_163 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_164 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15086) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_164 <= _pht_T_3;
        end else begin
          pht_7_164 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_165 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15089) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_165 <= _pht_T_3;
        end else begin
          pht_7_165 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_166 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15092) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_166 <= _pht_T_3;
        end else begin
          pht_7_166 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_167 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15095) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_167 <= _pht_T_3;
        end else begin
          pht_7_167 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_168 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15098) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_168 <= _pht_T_3;
        end else begin
          pht_7_168 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_169 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15101) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_169 <= _pht_T_3;
        end else begin
          pht_7_169 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_170 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15104) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_170 <= _pht_T_3;
        end else begin
          pht_7_170 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_171 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15107) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_171 <= _pht_T_3;
        end else begin
          pht_7_171 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_172 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15110) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_172 <= _pht_T_3;
        end else begin
          pht_7_172 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_173 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15113) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_173 <= _pht_T_3;
        end else begin
          pht_7_173 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_174 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15116) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_174 <= _pht_T_3;
        end else begin
          pht_7_174 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_175 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15119) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_175 <= _pht_T_3;
        end else begin
          pht_7_175 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_176 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15122) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_176 <= _pht_T_3;
        end else begin
          pht_7_176 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_177 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15125) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_177 <= _pht_T_3;
        end else begin
          pht_7_177 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_178 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15128) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_178 <= _pht_T_3;
        end else begin
          pht_7_178 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_179 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15131) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_179 <= _pht_T_3;
        end else begin
          pht_7_179 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_180 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15134) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_180 <= _pht_T_3;
        end else begin
          pht_7_180 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_181 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15137) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_181 <= _pht_T_3;
        end else begin
          pht_7_181 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_182 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15140) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_182 <= _pht_T_3;
        end else begin
          pht_7_182 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_183 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15143) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_183 <= _pht_T_3;
        end else begin
          pht_7_183 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_184 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15146) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_184 <= _pht_T_3;
        end else begin
          pht_7_184 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_185 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15149) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_185 <= _pht_T_3;
        end else begin
          pht_7_185 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_186 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15152) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_186 <= _pht_T_3;
        end else begin
          pht_7_186 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_187 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15155) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_187 <= _pht_T_3;
        end else begin
          pht_7_187 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_188 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15158) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_188 <= _pht_T_3;
        end else begin
          pht_7_188 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_189 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15161) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_189 <= _pht_T_3;
        end else begin
          pht_7_189 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_190 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15164) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_190 <= _pht_T_3;
        end else begin
          pht_7_190 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_191 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15167) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_191 <= _pht_T_3;
        end else begin
          pht_7_191 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_192 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15170) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_192 <= _pht_T_3;
        end else begin
          pht_7_192 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_193 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15173) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_193 <= _pht_T_3;
        end else begin
          pht_7_193 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_194 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15176) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_194 <= _pht_T_3;
        end else begin
          pht_7_194 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_195 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15179) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_195 <= _pht_T_3;
        end else begin
          pht_7_195 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_196 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15182) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_196 <= _pht_T_3;
        end else begin
          pht_7_196 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_197 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15185) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_197 <= _pht_T_3;
        end else begin
          pht_7_197 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_198 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15188) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_198 <= _pht_T_3;
        end else begin
          pht_7_198 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_199 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15191) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_199 <= _pht_T_3;
        end else begin
          pht_7_199 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_200 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15194) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_200 <= _pht_T_3;
        end else begin
          pht_7_200 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_201 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15197) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_201 <= _pht_T_3;
        end else begin
          pht_7_201 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_202 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15200) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_202 <= _pht_T_3;
        end else begin
          pht_7_202 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_203 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15203) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_203 <= _pht_T_3;
        end else begin
          pht_7_203 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_204 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15206) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_204 <= _pht_T_3;
        end else begin
          pht_7_204 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_205 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15209) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_205 <= _pht_T_3;
        end else begin
          pht_7_205 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_206 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15212) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_206 <= _pht_T_3;
        end else begin
          pht_7_206 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_207 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15215) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_207 <= _pht_T_3;
        end else begin
          pht_7_207 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_208 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15218) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_208 <= _pht_T_3;
        end else begin
          pht_7_208 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_209 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15221) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_209 <= _pht_T_3;
        end else begin
          pht_7_209 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_210 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15224) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_210 <= _pht_T_3;
        end else begin
          pht_7_210 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_211 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15227) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_211 <= _pht_T_3;
        end else begin
          pht_7_211 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_212 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15230) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_212 <= _pht_T_3;
        end else begin
          pht_7_212 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_213 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15233) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_213 <= _pht_T_3;
        end else begin
          pht_7_213 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_214 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15236) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_214 <= _pht_T_3;
        end else begin
          pht_7_214 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_215 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15239) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_215 <= _pht_T_3;
        end else begin
          pht_7_215 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_216 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15242) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_216 <= _pht_T_3;
        end else begin
          pht_7_216 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_217 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15245) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_217 <= _pht_T_3;
        end else begin
          pht_7_217 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_218 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15248) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_218 <= _pht_T_3;
        end else begin
          pht_7_218 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_219 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15251) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_219 <= _pht_T_3;
        end else begin
          pht_7_219 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_220 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15254) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_220 <= _pht_T_3;
        end else begin
          pht_7_220 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_221 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15257) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_221 <= _pht_T_3;
        end else begin
          pht_7_221 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_222 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15260) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_222 <= _pht_T_3;
        end else begin
          pht_7_222 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_223 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15263) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_223 <= _pht_T_3;
        end else begin
          pht_7_223 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_224 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15266) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_224 <= _pht_T_3;
        end else begin
          pht_7_224 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_225 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15269) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_225 <= _pht_T_3;
        end else begin
          pht_7_225 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_226 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15272) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_226 <= _pht_T_3;
        end else begin
          pht_7_226 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_227 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15275) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_227 <= _pht_T_3;
        end else begin
          pht_7_227 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_228 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15278) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_228 <= _pht_T_3;
        end else begin
          pht_7_228 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_229 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15281) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_229 <= _pht_T_3;
        end else begin
          pht_7_229 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_230 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15284) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_230 <= _pht_T_3;
        end else begin
          pht_7_230 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_231 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15287) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_231 <= _pht_T_3;
        end else begin
          pht_7_231 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_232 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15290) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_232 <= _pht_T_3;
        end else begin
          pht_7_232 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_233 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15293) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_233 <= _pht_T_3;
        end else begin
          pht_7_233 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_234 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15296) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_234 <= _pht_T_3;
        end else begin
          pht_7_234 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_235 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15299) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_235 <= _pht_T_3;
        end else begin
          pht_7_235 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_236 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15302) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_236 <= _pht_T_3;
        end else begin
          pht_7_236 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_237 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15305) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_237 <= _pht_T_3;
        end else begin
          pht_7_237 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_238 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15308) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_238 <= _pht_T_3;
        end else begin
          pht_7_238 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_239 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15311) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_239 <= _pht_T_3;
        end else begin
          pht_7_239 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_240 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15314) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_240 <= _pht_T_3;
        end else begin
          pht_7_240 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_241 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15317) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_241 <= _pht_T_3;
        end else begin
          pht_7_241 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_242 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15320) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_242 <= _pht_T_3;
        end else begin
          pht_7_242 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_243 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15323) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_243 <= _pht_T_3;
        end else begin
          pht_7_243 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_244 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15326) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_244 <= _pht_T_3;
        end else begin
          pht_7_244 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_245 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15329) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_245 <= _pht_T_3;
        end else begin
          pht_7_245 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_246 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15332) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_246 <= _pht_T_3;
        end else begin
          pht_7_246 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_247 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15335) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_247 <= _pht_T_3;
        end else begin
          pht_7_247 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_248 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15338) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_248 <= _pht_T_3;
        end else begin
          pht_7_248 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_249 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15341) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_249 <= _pht_T_3;
        end else begin
          pht_7_249 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_250 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15344) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_250 <= _pht_T_3;
        end else begin
          pht_7_250 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_251 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15347) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_251 <= _pht_T_3;
        end else begin
          pht_7_251 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_252 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15350) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_252 <= _pht_T_3;
        end else begin
          pht_7_252 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_253 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15353) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_253 <= _pht_T_3;
        end else begin
          pht_7_253 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_254 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15356) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_254 <= _pht_T_3;
        end else begin
          pht_7_254 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 51:20]
      pht_7_255 <= 2'h1; // @[BrPredictor.scala 51:20]
    end else if (io_jmp_packet_valid) begin // @[BrPredictor.scala 74:27]
      if (_GEN_19584 & _GEN_15359) begin // @[BrPredictor.scala 75:16]
        if (2'h3 == _GEN_4351) begin // @[Mux.scala 80:57]
          pht_7_255 <= _pht_T_3;
        end else begin
          pht_7_255 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_0_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_0_valid <= _GEN_8576;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_0_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h0 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_0_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_0_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h0 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_0_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_1_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_1_valid <= _GEN_8577;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_1_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_1_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_1_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_1_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_2_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_2_valid <= _GEN_8578;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_2_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_2_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_2_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_2_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_3_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_3_valid <= _GEN_8579;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_3_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_3_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_3_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_3_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_4_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_4_valid <= _GEN_8580;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_4_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h4 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_4_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_4_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h4 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_4_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_5_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_5_valid <= _GEN_8581;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_5_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h5 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_5_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_5_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h5 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_5_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_6_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_6_valid <= _GEN_8582;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_6_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h6 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_6_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_6_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h6 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_6_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_7_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_7_valid <= _GEN_8583;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_7_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h7 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_7_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_7_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h7 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_7_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_8_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_8_valid <= _GEN_8584;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_8_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h8 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_8_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_8_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h8 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_8_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_9_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_9_valid <= _GEN_8585;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_9_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h9 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_9_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_9_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h9 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_9_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_10_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_10_valid <= _GEN_8586;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_10_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'ha == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_10_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_10_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'ha == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_10_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_11_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_11_valid <= _GEN_8587;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_11_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'hb == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_11_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_11_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'hb == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_11_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_12_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_12_valid <= _GEN_8588;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_12_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'hc == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_12_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_12_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'hc == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_12_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_13_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_13_valid <= _GEN_8589;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_13_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'hd == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_13_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_13_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'hd == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_13_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_14_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_14_valid <= _GEN_8590;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_14_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'he == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_14_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_14_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'he == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_14_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_15_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_15_valid <= _GEN_8591;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_15_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'hf == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_15_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_15_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'hf == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_15_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_16_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_16_valid <= _GEN_8592;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_16_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h10 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_16_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_16_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h10 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_16_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_17_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_17_valid <= _GEN_8593;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_17_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h11 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_17_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_17_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h11 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_17_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_18_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_18_valid <= _GEN_8594;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_18_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h12 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_18_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_18_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h12 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_18_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_19_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_19_valid <= _GEN_8595;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_19_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h13 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_19_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_19_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h13 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_19_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_20_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_20_valid <= _GEN_8596;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_20_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h14 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_20_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_20_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h14 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_20_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_21_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_21_valid <= _GEN_8597;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_21_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h15 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_21_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_21_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h15 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_21_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_22_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_22_valid <= _GEN_8598;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_22_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h16 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_22_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_22_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h16 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_22_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_23_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_23_valid <= _GEN_8599;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_23_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h17 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_23_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_23_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h17 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_23_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_24_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_24_valid <= _GEN_8600;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_24_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h18 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_24_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_24_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h18 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_24_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_25_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_25_valid <= _GEN_8601;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_25_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h19 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_25_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_25_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h19 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_25_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_26_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_26_valid <= _GEN_8602;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_26_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1a == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_26_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_26_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1a == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_26_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_27_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_27_valid <= _GEN_8603;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_27_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1b == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_27_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_27_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1b == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_27_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_28_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_28_valid <= _GEN_8604;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_28_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1c == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_28_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_28_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1c == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_28_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_29_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_29_valid <= _GEN_8605;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_29_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1d == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_29_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_29_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1d == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_29_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_30_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_30_valid <= _GEN_8606;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_30_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1e == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_30_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_30_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1e == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_30_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_31_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_31_valid <= _GEN_8607;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_31_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1f == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_31_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_31_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h1f == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_31_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_32_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_32_valid <= _GEN_8608;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_32_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h20 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_32_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_32_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h20 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_32_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_33_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_33_valid <= _GEN_8609;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_33_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h21 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_33_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_33_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h21 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_33_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_34_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_34_valid <= _GEN_8610;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_34_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h22 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_34_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_34_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h22 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_34_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_35_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_35_valid <= _GEN_8611;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_35_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h23 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_35_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_35_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h23 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_35_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_36_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_36_valid <= _GEN_8612;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_36_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h24 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_36_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_36_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h24 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_36_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_37_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_37_valid <= _GEN_8613;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_37_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h25 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_37_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_37_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h25 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_37_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_38_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_38_valid <= _GEN_8614;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_38_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h26 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_38_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_38_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h26 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_38_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_39_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_39_valid <= _GEN_8615;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_39_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h27 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_39_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_39_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h27 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_39_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_40_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_40_valid <= _GEN_8616;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_40_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h28 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_40_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_40_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h28 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_40_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_41_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_41_valid <= _GEN_8617;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_41_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h29 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_41_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_41_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h29 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_41_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_42_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_42_valid <= _GEN_8618;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_42_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2a == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_42_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_42_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2a == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_42_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_43_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_43_valid <= _GEN_8619;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_43_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2b == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_43_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_43_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2b == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_43_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_44_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_44_valid <= _GEN_8620;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_44_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2c == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_44_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_44_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2c == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_44_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_45_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_45_valid <= _GEN_8621;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_45_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2d == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_45_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_45_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2d == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_45_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_46_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_46_valid <= _GEN_8622;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_46_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2e == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_46_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_46_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2e == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_46_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_47_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_47_valid <= _GEN_8623;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_47_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2f == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_47_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_47_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h2f == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_47_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_48_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_48_valid <= _GEN_8624;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_48_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h30 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_48_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_48_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h30 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_48_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_49_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_49_valid <= _GEN_8625;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_49_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h31 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_49_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_49_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h31 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_49_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_50_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_50_valid <= _GEN_8626;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_50_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h32 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_50_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_50_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h32 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_50_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_51_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_51_valid <= _GEN_8627;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_51_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h33 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_51_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_51_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h33 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_51_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_52_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_52_valid <= _GEN_8628;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_52_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h34 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_52_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_52_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h34 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_52_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_53_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_53_valid <= _GEN_8629;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_53_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h35 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_53_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_53_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h35 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_53_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_54_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_54_valid <= _GEN_8630;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_54_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h36 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_54_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_54_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h36 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_54_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_55_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_55_valid <= _GEN_8631;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_55_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h37 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_55_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_55_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h37 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_55_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_56_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_56_valid <= _GEN_8632;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_56_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h38 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_56_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_56_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h38 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_56_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_57_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_57_valid <= _GEN_8633;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_57_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h39 == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_57_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_57_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h39 == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_57_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_58_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_58_valid <= _GEN_8634;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_58_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3a == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_58_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_58_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3a == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_58_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_59_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_59_valid <= _GEN_8635;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_59_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3b == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_59_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_59_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3b == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_59_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_60_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_60_valid <= _GEN_8636;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_60_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3c == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_60_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_60_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3c == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_60_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_61_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_61_valid <= _GEN_8637;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_61_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3d == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_61_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_61_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3d == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_61_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_62_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_62_valid <= _GEN_8638;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_62_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3e == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_62_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_62_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3e == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_62_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_63_valid <= 1'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      btb_63_valid <= _GEN_8639;
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_63_tag <= 8'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3f == bht_waddr) begin // @[BrPredictor.scala 105:24]
        btb_63_tag <= io_jmp_packet_inst_pc[15:8]; // @[BrPredictor.scala 105:24]
      end
    end
    if (reset) begin // @[BrPredictor.scala 90:20]
      btb_63_target <= 32'h0; // @[BrPredictor.scala 90:20]
    end else if (io_jmp_packet_valid & io_jmp_packet_jmp) begin // @[BrPredictor.scala 103:45]
      if (6'h3f == bht_waddr) begin // @[BrPredictor.scala 106:27]
        btb_63_target <= io_jmp_packet_jmp_pc; // @[BrPredictor.scala 106:27]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bht_0 = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  bht_1 = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  bht_2 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  bht_3 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  bht_4 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  bht_5 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  bht_6 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  bht_7 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  bht_8 = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  bht_9 = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  bht_10 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  bht_11 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  bht_12 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  bht_13 = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  bht_14 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  bht_15 = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  bht_16 = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  bht_17 = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  bht_18 = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  bht_19 = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  bht_20 = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  bht_21 = _RAND_21[5:0];
  _RAND_22 = {1{`RANDOM}};
  bht_22 = _RAND_22[5:0];
  _RAND_23 = {1{`RANDOM}};
  bht_23 = _RAND_23[5:0];
  _RAND_24 = {1{`RANDOM}};
  bht_24 = _RAND_24[5:0];
  _RAND_25 = {1{`RANDOM}};
  bht_25 = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  bht_26 = _RAND_26[5:0];
  _RAND_27 = {1{`RANDOM}};
  bht_27 = _RAND_27[5:0];
  _RAND_28 = {1{`RANDOM}};
  bht_28 = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  bht_29 = _RAND_29[5:0];
  _RAND_30 = {1{`RANDOM}};
  bht_30 = _RAND_30[5:0];
  _RAND_31 = {1{`RANDOM}};
  bht_31 = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  bht_32 = _RAND_32[5:0];
  _RAND_33 = {1{`RANDOM}};
  bht_33 = _RAND_33[5:0];
  _RAND_34 = {1{`RANDOM}};
  bht_34 = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  bht_35 = _RAND_35[5:0];
  _RAND_36 = {1{`RANDOM}};
  bht_36 = _RAND_36[5:0];
  _RAND_37 = {1{`RANDOM}};
  bht_37 = _RAND_37[5:0];
  _RAND_38 = {1{`RANDOM}};
  bht_38 = _RAND_38[5:0];
  _RAND_39 = {1{`RANDOM}};
  bht_39 = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
  bht_40 = _RAND_40[5:0];
  _RAND_41 = {1{`RANDOM}};
  bht_41 = _RAND_41[5:0];
  _RAND_42 = {1{`RANDOM}};
  bht_42 = _RAND_42[5:0];
  _RAND_43 = {1{`RANDOM}};
  bht_43 = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  bht_44 = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  bht_45 = _RAND_45[5:0];
  _RAND_46 = {1{`RANDOM}};
  bht_46 = _RAND_46[5:0];
  _RAND_47 = {1{`RANDOM}};
  bht_47 = _RAND_47[5:0];
  _RAND_48 = {1{`RANDOM}};
  bht_48 = _RAND_48[5:0];
  _RAND_49 = {1{`RANDOM}};
  bht_49 = _RAND_49[5:0];
  _RAND_50 = {1{`RANDOM}};
  bht_50 = _RAND_50[5:0];
  _RAND_51 = {1{`RANDOM}};
  bht_51 = _RAND_51[5:0];
  _RAND_52 = {1{`RANDOM}};
  bht_52 = _RAND_52[5:0];
  _RAND_53 = {1{`RANDOM}};
  bht_53 = _RAND_53[5:0];
  _RAND_54 = {1{`RANDOM}};
  bht_54 = _RAND_54[5:0];
  _RAND_55 = {1{`RANDOM}};
  bht_55 = _RAND_55[5:0];
  _RAND_56 = {1{`RANDOM}};
  bht_56 = _RAND_56[5:0];
  _RAND_57 = {1{`RANDOM}};
  bht_57 = _RAND_57[5:0];
  _RAND_58 = {1{`RANDOM}};
  bht_58 = _RAND_58[5:0];
  _RAND_59 = {1{`RANDOM}};
  bht_59 = _RAND_59[5:0];
  _RAND_60 = {1{`RANDOM}};
  bht_60 = _RAND_60[5:0];
  _RAND_61 = {1{`RANDOM}};
  bht_61 = _RAND_61[5:0];
  _RAND_62 = {1{`RANDOM}};
  bht_62 = _RAND_62[5:0];
  _RAND_63 = {1{`RANDOM}};
  bht_63 = _RAND_63[5:0];
  _RAND_64 = {1{`RANDOM}};
  pht_0_0 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  pht_0_1 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  pht_0_2 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  pht_0_3 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  pht_0_4 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  pht_0_5 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  pht_0_6 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  pht_0_7 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  pht_0_8 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  pht_0_9 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  pht_0_10 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  pht_0_11 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  pht_0_12 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  pht_0_13 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  pht_0_14 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  pht_0_15 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  pht_0_16 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  pht_0_17 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  pht_0_18 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  pht_0_19 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  pht_0_20 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  pht_0_21 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  pht_0_22 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  pht_0_23 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  pht_0_24 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  pht_0_25 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  pht_0_26 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  pht_0_27 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  pht_0_28 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  pht_0_29 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  pht_0_30 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  pht_0_31 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  pht_0_32 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  pht_0_33 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  pht_0_34 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  pht_0_35 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  pht_0_36 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  pht_0_37 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  pht_0_38 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  pht_0_39 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  pht_0_40 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  pht_0_41 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  pht_0_42 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  pht_0_43 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  pht_0_44 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  pht_0_45 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  pht_0_46 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  pht_0_47 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  pht_0_48 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  pht_0_49 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  pht_0_50 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  pht_0_51 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  pht_0_52 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  pht_0_53 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  pht_0_54 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  pht_0_55 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  pht_0_56 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  pht_0_57 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  pht_0_58 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  pht_0_59 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  pht_0_60 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  pht_0_61 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  pht_0_62 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  pht_0_63 = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  pht_0_64 = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  pht_0_65 = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  pht_0_66 = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  pht_0_67 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  pht_0_68 = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  pht_0_69 = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  pht_0_70 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  pht_0_71 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  pht_0_72 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  pht_0_73 = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  pht_0_74 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  pht_0_75 = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  pht_0_76 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  pht_0_77 = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  pht_0_78 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  pht_0_79 = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  pht_0_80 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  pht_0_81 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  pht_0_82 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  pht_0_83 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  pht_0_84 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  pht_0_85 = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  pht_0_86 = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  pht_0_87 = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  pht_0_88 = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  pht_0_89 = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  pht_0_90 = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  pht_0_91 = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  pht_0_92 = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  pht_0_93 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  pht_0_94 = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  pht_0_95 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  pht_0_96 = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  pht_0_97 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  pht_0_98 = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  pht_0_99 = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  pht_0_100 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  pht_0_101 = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  pht_0_102 = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  pht_0_103 = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  pht_0_104 = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  pht_0_105 = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  pht_0_106 = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  pht_0_107 = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  pht_0_108 = _RAND_172[1:0];
  _RAND_173 = {1{`RANDOM}};
  pht_0_109 = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  pht_0_110 = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  pht_0_111 = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  pht_0_112 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  pht_0_113 = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  pht_0_114 = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  pht_0_115 = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  pht_0_116 = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  pht_0_117 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  pht_0_118 = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  pht_0_119 = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  pht_0_120 = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  pht_0_121 = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  pht_0_122 = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  pht_0_123 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  pht_0_124 = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  pht_0_125 = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  pht_0_126 = _RAND_190[1:0];
  _RAND_191 = {1{`RANDOM}};
  pht_0_127 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  pht_0_128 = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  pht_0_129 = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  pht_0_130 = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  pht_0_131 = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  pht_0_132 = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  pht_0_133 = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  pht_0_134 = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  pht_0_135 = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  pht_0_136 = _RAND_200[1:0];
  _RAND_201 = {1{`RANDOM}};
  pht_0_137 = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  pht_0_138 = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  pht_0_139 = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  pht_0_140 = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  pht_0_141 = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  pht_0_142 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  pht_0_143 = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  pht_0_144 = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  pht_0_145 = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  pht_0_146 = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  pht_0_147 = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  pht_0_148 = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  pht_0_149 = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  pht_0_150 = _RAND_214[1:0];
  _RAND_215 = {1{`RANDOM}};
  pht_0_151 = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  pht_0_152 = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  pht_0_153 = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  pht_0_154 = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  pht_0_155 = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  pht_0_156 = _RAND_220[1:0];
  _RAND_221 = {1{`RANDOM}};
  pht_0_157 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  pht_0_158 = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  pht_0_159 = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  pht_0_160 = _RAND_224[1:0];
  _RAND_225 = {1{`RANDOM}};
  pht_0_161 = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  pht_0_162 = _RAND_226[1:0];
  _RAND_227 = {1{`RANDOM}};
  pht_0_163 = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  pht_0_164 = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  pht_0_165 = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  pht_0_166 = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  pht_0_167 = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  pht_0_168 = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  pht_0_169 = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  pht_0_170 = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  pht_0_171 = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  pht_0_172 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  pht_0_173 = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  pht_0_174 = _RAND_238[1:0];
  _RAND_239 = {1{`RANDOM}};
  pht_0_175 = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  pht_0_176 = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  pht_0_177 = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  pht_0_178 = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  pht_0_179 = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  pht_0_180 = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  pht_0_181 = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  pht_0_182 = _RAND_246[1:0];
  _RAND_247 = {1{`RANDOM}};
  pht_0_183 = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  pht_0_184 = _RAND_248[1:0];
  _RAND_249 = {1{`RANDOM}};
  pht_0_185 = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  pht_0_186 = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  pht_0_187 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  pht_0_188 = _RAND_252[1:0];
  _RAND_253 = {1{`RANDOM}};
  pht_0_189 = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  pht_0_190 = _RAND_254[1:0];
  _RAND_255 = {1{`RANDOM}};
  pht_0_191 = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  pht_0_192 = _RAND_256[1:0];
  _RAND_257 = {1{`RANDOM}};
  pht_0_193 = _RAND_257[1:0];
  _RAND_258 = {1{`RANDOM}};
  pht_0_194 = _RAND_258[1:0];
  _RAND_259 = {1{`RANDOM}};
  pht_0_195 = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  pht_0_196 = _RAND_260[1:0];
  _RAND_261 = {1{`RANDOM}};
  pht_0_197 = _RAND_261[1:0];
  _RAND_262 = {1{`RANDOM}};
  pht_0_198 = _RAND_262[1:0];
  _RAND_263 = {1{`RANDOM}};
  pht_0_199 = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  pht_0_200 = _RAND_264[1:0];
  _RAND_265 = {1{`RANDOM}};
  pht_0_201 = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  pht_0_202 = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  pht_0_203 = _RAND_267[1:0];
  _RAND_268 = {1{`RANDOM}};
  pht_0_204 = _RAND_268[1:0];
  _RAND_269 = {1{`RANDOM}};
  pht_0_205 = _RAND_269[1:0];
  _RAND_270 = {1{`RANDOM}};
  pht_0_206 = _RAND_270[1:0];
  _RAND_271 = {1{`RANDOM}};
  pht_0_207 = _RAND_271[1:0];
  _RAND_272 = {1{`RANDOM}};
  pht_0_208 = _RAND_272[1:0];
  _RAND_273 = {1{`RANDOM}};
  pht_0_209 = _RAND_273[1:0];
  _RAND_274 = {1{`RANDOM}};
  pht_0_210 = _RAND_274[1:0];
  _RAND_275 = {1{`RANDOM}};
  pht_0_211 = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  pht_0_212 = _RAND_276[1:0];
  _RAND_277 = {1{`RANDOM}};
  pht_0_213 = _RAND_277[1:0];
  _RAND_278 = {1{`RANDOM}};
  pht_0_214 = _RAND_278[1:0];
  _RAND_279 = {1{`RANDOM}};
  pht_0_215 = _RAND_279[1:0];
  _RAND_280 = {1{`RANDOM}};
  pht_0_216 = _RAND_280[1:0];
  _RAND_281 = {1{`RANDOM}};
  pht_0_217 = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  pht_0_218 = _RAND_282[1:0];
  _RAND_283 = {1{`RANDOM}};
  pht_0_219 = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  pht_0_220 = _RAND_284[1:0];
  _RAND_285 = {1{`RANDOM}};
  pht_0_221 = _RAND_285[1:0];
  _RAND_286 = {1{`RANDOM}};
  pht_0_222 = _RAND_286[1:0];
  _RAND_287 = {1{`RANDOM}};
  pht_0_223 = _RAND_287[1:0];
  _RAND_288 = {1{`RANDOM}};
  pht_0_224 = _RAND_288[1:0];
  _RAND_289 = {1{`RANDOM}};
  pht_0_225 = _RAND_289[1:0];
  _RAND_290 = {1{`RANDOM}};
  pht_0_226 = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  pht_0_227 = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  pht_0_228 = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  pht_0_229 = _RAND_293[1:0];
  _RAND_294 = {1{`RANDOM}};
  pht_0_230 = _RAND_294[1:0];
  _RAND_295 = {1{`RANDOM}};
  pht_0_231 = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  pht_0_232 = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  pht_0_233 = _RAND_297[1:0];
  _RAND_298 = {1{`RANDOM}};
  pht_0_234 = _RAND_298[1:0];
  _RAND_299 = {1{`RANDOM}};
  pht_0_235 = _RAND_299[1:0];
  _RAND_300 = {1{`RANDOM}};
  pht_0_236 = _RAND_300[1:0];
  _RAND_301 = {1{`RANDOM}};
  pht_0_237 = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  pht_0_238 = _RAND_302[1:0];
  _RAND_303 = {1{`RANDOM}};
  pht_0_239 = _RAND_303[1:0];
  _RAND_304 = {1{`RANDOM}};
  pht_0_240 = _RAND_304[1:0];
  _RAND_305 = {1{`RANDOM}};
  pht_0_241 = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  pht_0_242 = _RAND_306[1:0];
  _RAND_307 = {1{`RANDOM}};
  pht_0_243 = _RAND_307[1:0];
  _RAND_308 = {1{`RANDOM}};
  pht_0_244 = _RAND_308[1:0];
  _RAND_309 = {1{`RANDOM}};
  pht_0_245 = _RAND_309[1:0];
  _RAND_310 = {1{`RANDOM}};
  pht_0_246 = _RAND_310[1:0];
  _RAND_311 = {1{`RANDOM}};
  pht_0_247 = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  pht_0_248 = _RAND_312[1:0];
  _RAND_313 = {1{`RANDOM}};
  pht_0_249 = _RAND_313[1:0];
  _RAND_314 = {1{`RANDOM}};
  pht_0_250 = _RAND_314[1:0];
  _RAND_315 = {1{`RANDOM}};
  pht_0_251 = _RAND_315[1:0];
  _RAND_316 = {1{`RANDOM}};
  pht_0_252 = _RAND_316[1:0];
  _RAND_317 = {1{`RANDOM}};
  pht_0_253 = _RAND_317[1:0];
  _RAND_318 = {1{`RANDOM}};
  pht_0_254 = _RAND_318[1:0];
  _RAND_319 = {1{`RANDOM}};
  pht_0_255 = _RAND_319[1:0];
  _RAND_320 = {1{`RANDOM}};
  pht_1_0 = _RAND_320[1:0];
  _RAND_321 = {1{`RANDOM}};
  pht_1_1 = _RAND_321[1:0];
  _RAND_322 = {1{`RANDOM}};
  pht_1_2 = _RAND_322[1:0];
  _RAND_323 = {1{`RANDOM}};
  pht_1_3 = _RAND_323[1:0];
  _RAND_324 = {1{`RANDOM}};
  pht_1_4 = _RAND_324[1:0];
  _RAND_325 = {1{`RANDOM}};
  pht_1_5 = _RAND_325[1:0];
  _RAND_326 = {1{`RANDOM}};
  pht_1_6 = _RAND_326[1:0];
  _RAND_327 = {1{`RANDOM}};
  pht_1_7 = _RAND_327[1:0];
  _RAND_328 = {1{`RANDOM}};
  pht_1_8 = _RAND_328[1:0];
  _RAND_329 = {1{`RANDOM}};
  pht_1_9 = _RAND_329[1:0];
  _RAND_330 = {1{`RANDOM}};
  pht_1_10 = _RAND_330[1:0];
  _RAND_331 = {1{`RANDOM}};
  pht_1_11 = _RAND_331[1:0];
  _RAND_332 = {1{`RANDOM}};
  pht_1_12 = _RAND_332[1:0];
  _RAND_333 = {1{`RANDOM}};
  pht_1_13 = _RAND_333[1:0];
  _RAND_334 = {1{`RANDOM}};
  pht_1_14 = _RAND_334[1:0];
  _RAND_335 = {1{`RANDOM}};
  pht_1_15 = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  pht_1_16 = _RAND_336[1:0];
  _RAND_337 = {1{`RANDOM}};
  pht_1_17 = _RAND_337[1:0];
  _RAND_338 = {1{`RANDOM}};
  pht_1_18 = _RAND_338[1:0];
  _RAND_339 = {1{`RANDOM}};
  pht_1_19 = _RAND_339[1:0];
  _RAND_340 = {1{`RANDOM}};
  pht_1_20 = _RAND_340[1:0];
  _RAND_341 = {1{`RANDOM}};
  pht_1_21 = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  pht_1_22 = _RAND_342[1:0];
  _RAND_343 = {1{`RANDOM}};
  pht_1_23 = _RAND_343[1:0];
  _RAND_344 = {1{`RANDOM}};
  pht_1_24 = _RAND_344[1:0];
  _RAND_345 = {1{`RANDOM}};
  pht_1_25 = _RAND_345[1:0];
  _RAND_346 = {1{`RANDOM}};
  pht_1_26 = _RAND_346[1:0];
  _RAND_347 = {1{`RANDOM}};
  pht_1_27 = _RAND_347[1:0];
  _RAND_348 = {1{`RANDOM}};
  pht_1_28 = _RAND_348[1:0];
  _RAND_349 = {1{`RANDOM}};
  pht_1_29 = _RAND_349[1:0];
  _RAND_350 = {1{`RANDOM}};
  pht_1_30 = _RAND_350[1:0];
  _RAND_351 = {1{`RANDOM}};
  pht_1_31 = _RAND_351[1:0];
  _RAND_352 = {1{`RANDOM}};
  pht_1_32 = _RAND_352[1:0];
  _RAND_353 = {1{`RANDOM}};
  pht_1_33 = _RAND_353[1:0];
  _RAND_354 = {1{`RANDOM}};
  pht_1_34 = _RAND_354[1:0];
  _RAND_355 = {1{`RANDOM}};
  pht_1_35 = _RAND_355[1:0];
  _RAND_356 = {1{`RANDOM}};
  pht_1_36 = _RAND_356[1:0];
  _RAND_357 = {1{`RANDOM}};
  pht_1_37 = _RAND_357[1:0];
  _RAND_358 = {1{`RANDOM}};
  pht_1_38 = _RAND_358[1:0];
  _RAND_359 = {1{`RANDOM}};
  pht_1_39 = _RAND_359[1:0];
  _RAND_360 = {1{`RANDOM}};
  pht_1_40 = _RAND_360[1:0];
  _RAND_361 = {1{`RANDOM}};
  pht_1_41 = _RAND_361[1:0];
  _RAND_362 = {1{`RANDOM}};
  pht_1_42 = _RAND_362[1:0];
  _RAND_363 = {1{`RANDOM}};
  pht_1_43 = _RAND_363[1:0];
  _RAND_364 = {1{`RANDOM}};
  pht_1_44 = _RAND_364[1:0];
  _RAND_365 = {1{`RANDOM}};
  pht_1_45 = _RAND_365[1:0];
  _RAND_366 = {1{`RANDOM}};
  pht_1_46 = _RAND_366[1:0];
  _RAND_367 = {1{`RANDOM}};
  pht_1_47 = _RAND_367[1:0];
  _RAND_368 = {1{`RANDOM}};
  pht_1_48 = _RAND_368[1:0];
  _RAND_369 = {1{`RANDOM}};
  pht_1_49 = _RAND_369[1:0];
  _RAND_370 = {1{`RANDOM}};
  pht_1_50 = _RAND_370[1:0];
  _RAND_371 = {1{`RANDOM}};
  pht_1_51 = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  pht_1_52 = _RAND_372[1:0];
  _RAND_373 = {1{`RANDOM}};
  pht_1_53 = _RAND_373[1:0];
  _RAND_374 = {1{`RANDOM}};
  pht_1_54 = _RAND_374[1:0];
  _RAND_375 = {1{`RANDOM}};
  pht_1_55 = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  pht_1_56 = _RAND_376[1:0];
  _RAND_377 = {1{`RANDOM}};
  pht_1_57 = _RAND_377[1:0];
  _RAND_378 = {1{`RANDOM}};
  pht_1_58 = _RAND_378[1:0];
  _RAND_379 = {1{`RANDOM}};
  pht_1_59 = _RAND_379[1:0];
  _RAND_380 = {1{`RANDOM}};
  pht_1_60 = _RAND_380[1:0];
  _RAND_381 = {1{`RANDOM}};
  pht_1_61 = _RAND_381[1:0];
  _RAND_382 = {1{`RANDOM}};
  pht_1_62 = _RAND_382[1:0];
  _RAND_383 = {1{`RANDOM}};
  pht_1_63 = _RAND_383[1:0];
  _RAND_384 = {1{`RANDOM}};
  pht_1_64 = _RAND_384[1:0];
  _RAND_385 = {1{`RANDOM}};
  pht_1_65 = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  pht_1_66 = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  pht_1_67 = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  pht_1_68 = _RAND_388[1:0];
  _RAND_389 = {1{`RANDOM}};
  pht_1_69 = _RAND_389[1:0];
  _RAND_390 = {1{`RANDOM}};
  pht_1_70 = _RAND_390[1:0];
  _RAND_391 = {1{`RANDOM}};
  pht_1_71 = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  pht_1_72 = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  pht_1_73 = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  pht_1_74 = _RAND_394[1:0];
  _RAND_395 = {1{`RANDOM}};
  pht_1_75 = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  pht_1_76 = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  pht_1_77 = _RAND_397[1:0];
  _RAND_398 = {1{`RANDOM}};
  pht_1_78 = _RAND_398[1:0];
  _RAND_399 = {1{`RANDOM}};
  pht_1_79 = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  pht_1_80 = _RAND_400[1:0];
  _RAND_401 = {1{`RANDOM}};
  pht_1_81 = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  pht_1_82 = _RAND_402[1:0];
  _RAND_403 = {1{`RANDOM}};
  pht_1_83 = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  pht_1_84 = _RAND_404[1:0];
  _RAND_405 = {1{`RANDOM}};
  pht_1_85 = _RAND_405[1:0];
  _RAND_406 = {1{`RANDOM}};
  pht_1_86 = _RAND_406[1:0];
  _RAND_407 = {1{`RANDOM}};
  pht_1_87 = _RAND_407[1:0];
  _RAND_408 = {1{`RANDOM}};
  pht_1_88 = _RAND_408[1:0];
  _RAND_409 = {1{`RANDOM}};
  pht_1_89 = _RAND_409[1:0];
  _RAND_410 = {1{`RANDOM}};
  pht_1_90 = _RAND_410[1:0];
  _RAND_411 = {1{`RANDOM}};
  pht_1_91 = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  pht_1_92 = _RAND_412[1:0];
  _RAND_413 = {1{`RANDOM}};
  pht_1_93 = _RAND_413[1:0];
  _RAND_414 = {1{`RANDOM}};
  pht_1_94 = _RAND_414[1:0];
  _RAND_415 = {1{`RANDOM}};
  pht_1_95 = _RAND_415[1:0];
  _RAND_416 = {1{`RANDOM}};
  pht_1_96 = _RAND_416[1:0];
  _RAND_417 = {1{`RANDOM}};
  pht_1_97 = _RAND_417[1:0];
  _RAND_418 = {1{`RANDOM}};
  pht_1_98 = _RAND_418[1:0];
  _RAND_419 = {1{`RANDOM}};
  pht_1_99 = _RAND_419[1:0];
  _RAND_420 = {1{`RANDOM}};
  pht_1_100 = _RAND_420[1:0];
  _RAND_421 = {1{`RANDOM}};
  pht_1_101 = _RAND_421[1:0];
  _RAND_422 = {1{`RANDOM}};
  pht_1_102 = _RAND_422[1:0];
  _RAND_423 = {1{`RANDOM}};
  pht_1_103 = _RAND_423[1:0];
  _RAND_424 = {1{`RANDOM}};
  pht_1_104 = _RAND_424[1:0];
  _RAND_425 = {1{`RANDOM}};
  pht_1_105 = _RAND_425[1:0];
  _RAND_426 = {1{`RANDOM}};
  pht_1_106 = _RAND_426[1:0];
  _RAND_427 = {1{`RANDOM}};
  pht_1_107 = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  pht_1_108 = _RAND_428[1:0];
  _RAND_429 = {1{`RANDOM}};
  pht_1_109 = _RAND_429[1:0];
  _RAND_430 = {1{`RANDOM}};
  pht_1_110 = _RAND_430[1:0];
  _RAND_431 = {1{`RANDOM}};
  pht_1_111 = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  pht_1_112 = _RAND_432[1:0];
  _RAND_433 = {1{`RANDOM}};
  pht_1_113 = _RAND_433[1:0];
  _RAND_434 = {1{`RANDOM}};
  pht_1_114 = _RAND_434[1:0];
  _RAND_435 = {1{`RANDOM}};
  pht_1_115 = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  pht_1_116 = _RAND_436[1:0];
  _RAND_437 = {1{`RANDOM}};
  pht_1_117 = _RAND_437[1:0];
  _RAND_438 = {1{`RANDOM}};
  pht_1_118 = _RAND_438[1:0];
  _RAND_439 = {1{`RANDOM}};
  pht_1_119 = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  pht_1_120 = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  pht_1_121 = _RAND_441[1:0];
  _RAND_442 = {1{`RANDOM}};
  pht_1_122 = _RAND_442[1:0];
  _RAND_443 = {1{`RANDOM}};
  pht_1_123 = _RAND_443[1:0];
  _RAND_444 = {1{`RANDOM}};
  pht_1_124 = _RAND_444[1:0];
  _RAND_445 = {1{`RANDOM}};
  pht_1_125 = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  pht_1_126 = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  pht_1_127 = _RAND_447[1:0];
  _RAND_448 = {1{`RANDOM}};
  pht_1_128 = _RAND_448[1:0];
  _RAND_449 = {1{`RANDOM}};
  pht_1_129 = _RAND_449[1:0];
  _RAND_450 = {1{`RANDOM}};
  pht_1_130 = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  pht_1_131 = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  pht_1_132 = _RAND_452[1:0];
  _RAND_453 = {1{`RANDOM}};
  pht_1_133 = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  pht_1_134 = _RAND_454[1:0];
  _RAND_455 = {1{`RANDOM}};
  pht_1_135 = _RAND_455[1:0];
  _RAND_456 = {1{`RANDOM}};
  pht_1_136 = _RAND_456[1:0];
  _RAND_457 = {1{`RANDOM}};
  pht_1_137 = _RAND_457[1:0];
  _RAND_458 = {1{`RANDOM}};
  pht_1_138 = _RAND_458[1:0];
  _RAND_459 = {1{`RANDOM}};
  pht_1_139 = _RAND_459[1:0];
  _RAND_460 = {1{`RANDOM}};
  pht_1_140 = _RAND_460[1:0];
  _RAND_461 = {1{`RANDOM}};
  pht_1_141 = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  pht_1_142 = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  pht_1_143 = _RAND_463[1:0];
  _RAND_464 = {1{`RANDOM}};
  pht_1_144 = _RAND_464[1:0];
  _RAND_465 = {1{`RANDOM}};
  pht_1_145 = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  pht_1_146 = _RAND_466[1:0];
  _RAND_467 = {1{`RANDOM}};
  pht_1_147 = _RAND_467[1:0];
  _RAND_468 = {1{`RANDOM}};
  pht_1_148 = _RAND_468[1:0];
  _RAND_469 = {1{`RANDOM}};
  pht_1_149 = _RAND_469[1:0];
  _RAND_470 = {1{`RANDOM}};
  pht_1_150 = _RAND_470[1:0];
  _RAND_471 = {1{`RANDOM}};
  pht_1_151 = _RAND_471[1:0];
  _RAND_472 = {1{`RANDOM}};
  pht_1_152 = _RAND_472[1:0];
  _RAND_473 = {1{`RANDOM}};
  pht_1_153 = _RAND_473[1:0];
  _RAND_474 = {1{`RANDOM}};
  pht_1_154 = _RAND_474[1:0];
  _RAND_475 = {1{`RANDOM}};
  pht_1_155 = _RAND_475[1:0];
  _RAND_476 = {1{`RANDOM}};
  pht_1_156 = _RAND_476[1:0];
  _RAND_477 = {1{`RANDOM}};
  pht_1_157 = _RAND_477[1:0];
  _RAND_478 = {1{`RANDOM}};
  pht_1_158 = _RAND_478[1:0];
  _RAND_479 = {1{`RANDOM}};
  pht_1_159 = _RAND_479[1:0];
  _RAND_480 = {1{`RANDOM}};
  pht_1_160 = _RAND_480[1:0];
  _RAND_481 = {1{`RANDOM}};
  pht_1_161 = _RAND_481[1:0];
  _RAND_482 = {1{`RANDOM}};
  pht_1_162 = _RAND_482[1:0];
  _RAND_483 = {1{`RANDOM}};
  pht_1_163 = _RAND_483[1:0];
  _RAND_484 = {1{`RANDOM}};
  pht_1_164 = _RAND_484[1:0];
  _RAND_485 = {1{`RANDOM}};
  pht_1_165 = _RAND_485[1:0];
  _RAND_486 = {1{`RANDOM}};
  pht_1_166 = _RAND_486[1:0];
  _RAND_487 = {1{`RANDOM}};
  pht_1_167 = _RAND_487[1:0];
  _RAND_488 = {1{`RANDOM}};
  pht_1_168 = _RAND_488[1:0];
  _RAND_489 = {1{`RANDOM}};
  pht_1_169 = _RAND_489[1:0];
  _RAND_490 = {1{`RANDOM}};
  pht_1_170 = _RAND_490[1:0];
  _RAND_491 = {1{`RANDOM}};
  pht_1_171 = _RAND_491[1:0];
  _RAND_492 = {1{`RANDOM}};
  pht_1_172 = _RAND_492[1:0];
  _RAND_493 = {1{`RANDOM}};
  pht_1_173 = _RAND_493[1:0];
  _RAND_494 = {1{`RANDOM}};
  pht_1_174 = _RAND_494[1:0];
  _RAND_495 = {1{`RANDOM}};
  pht_1_175 = _RAND_495[1:0];
  _RAND_496 = {1{`RANDOM}};
  pht_1_176 = _RAND_496[1:0];
  _RAND_497 = {1{`RANDOM}};
  pht_1_177 = _RAND_497[1:0];
  _RAND_498 = {1{`RANDOM}};
  pht_1_178 = _RAND_498[1:0];
  _RAND_499 = {1{`RANDOM}};
  pht_1_179 = _RAND_499[1:0];
  _RAND_500 = {1{`RANDOM}};
  pht_1_180 = _RAND_500[1:0];
  _RAND_501 = {1{`RANDOM}};
  pht_1_181 = _RAND_501[1:0];
  _RAND_502 = {1{`RANDOM}};
  pht_1_182 = _RAND_502[1:0];
  _RAND_503 = {1{`RANDOM}};
  pht_1_183 = _RAND_503[1:0];
  _RAND_504 = {1{`RANDOM}};
  pht_1_184 = _RAND_504[1:0];
  _RAND_505 = {1{`RANDOM}};
  pht_1_185 = _RAND_505[1:0];
  _RAND_506 = {1{`RANDOM}};
  pht_1_186 = _RAND_506[1:0];
  _RAND_507 = {1{`RANDOM}};
  pht_1_187 = _RAND_507[1:0];
  _RAND_508 = {1{`RANDOM}};
  pht_1_188 = _RAND_508[1:0];
  _RAND_509 = {1{`RANDOM}};
  pht_1_189 = _RAND_509[1:0];
  _RAND_510 = {1{`RANDOM}};
  pht_1_190 = _RAND_510[1:0];
  _RAND_511 = {1{`RANDOM}};
  pht_1_191 = _RAND_511[1:0];
  _RAND_512 = {1{`RANDOM}};
  pht_1_192 = _RAND_512[1:0];
  _RAND_513 = {1{`RANDOM}};
  pht_1_193 = _RAND_513[1:0];
  _RAND_514 = {1{`RANDOM}};
  pht_1_194 = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  pht_1_195 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  pht_1_196 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  pht_1_197 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  pht_1_198 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  pht_1_199 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  pht_1_200 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  pht_1_201 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  pht_1_202 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  pht_1_203 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  pht_1_204 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  pht_1_205 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  pht_1_206 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  pht_1_207 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  pht_1_208 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  pht_1_209 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  pht_1_210 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  pht_1_211 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  pht_1_212 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  pht_1_213 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  pht_1_214 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  pht_1_215 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  pht_1_216 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  pht_1_217 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  pht_1_218 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  pht_1_219 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  pht_1_220 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  pht_1_221 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  pht_1_222 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  pht_1_223 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  pht_1_224 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  pht_1_225 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  pht_1_226 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  pht_1_227 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  pht_1_228 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  pht_1_229 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  pht_1_230 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  pht_1_231 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  pht_1_232 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  pht_1_233 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  pht_1_234 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  pht_1_235 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  pht_1_236 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  pht_1_237 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  pht_1_238 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  pht_1_239 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  pht_1_240 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  pht_1_241 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  pht_1_242 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  pht_1_243 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  pht_1_244 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  pht_1_245 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  pht_1_246 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  pht_1_247 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  pht_1_248 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  pht_1_249 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  pht_1_250 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  pht_1_251 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  pht_1_252 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  pht_1_253 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  pht_1_254 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  pht_1_255 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  pht_2_0 = _RAND_576[1:0];
  _RAND_577 = {1{`RANDOM}};
  pht_2_1 = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  pht_2_2 = _RAND_578[1:0];
  _RAND_579 = {1{`RANDOM}};
  pht_2_3 = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  pht_2_4 = _RAND_580[1:0];
  _RAND_581 = {1{`RANDOM}};
  pht_2_5 = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  pht_2_6 = _RAND_582[1:0];
  _RAND_583 = {1{`RANDOM}};
  pht_2_7 = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  pht_2_8 = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  pht_2_9 = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  pht_2_10 = _RAND_586[1:0];
  _RAND_587 = {1{`RANDOM}};
  pht_2_11 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  pht_2_12 = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  pht_2_13 = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  pht_2_14 = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  pht_2_15 = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  pht_2_16 = _RAND_592[1:0];
  _RAND_593 = {1{`RANDOM}};
  pht_2_17 = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  pht_2_18 = _RAND_594[1:0];
  _RAND_595 = {1{`RANDOM}};
  pht_2_19 = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  pht_2_20 = _RAND_596[1:0];
  _RAND_597 = {1{`RANDOM}};
  pht_2_21 = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  pht_2_22 = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  pht_2_23 = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  pht_2_24 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  pht_2_25 = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  pht_2_26 = _RAND_602[1:0];
  _RAND_603 = {1{`RANDOM}};
  pht_2_27 = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  pht_2_28 = _RAND_604[1:0];
  _RAND_605 = {1{`RANDOM}};
  pht_2_29 = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  pht_2_30 = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  pht_2_31 = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  pht_2_32 = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  pht_2_33 = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  pht_2_34 = _RAND_610[1:0];
  _RAND_611 = {1{`RANDOM}};
  pht_2_35 = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  pht_2_36 = _RAND_612[1:0];
  _RAND_613 = {1{`RANDOM}};
  pht_2_37 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  pht_2_38 = _RAND_614[1:0];
  _RAND_615 = {1{`RANDOM}};
  pht_2_39 = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  pht_2_40 = _RAND_616[1:0];
  _RAND_617 = {1{`RANDOM}};
  pht_2_41 = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  pht_2_42 = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  pht_2_43 = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  pht_2_44 = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  pht_2_45 = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  pht_2_46 = _RAND_622[1:0];
  _RAND_623 = {1{`RANDOM}};
  pht_2_47 = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  pht_2_48 = _RAND_624[1:0];
  _RAND_625 = {1{`RANDOM}};
  pht_2_49 = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  pht_2_50 = _RAND_626[1:0];
  _RAND_627 = {1{`RANDOM}};
  pht_2_51 = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  pht_2_52 = _RAND_628[1:0];
  _RAND_629 = {1{`RANDOM}};
  pht_2_53 = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  pht_2_54 = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  pht_2_55 = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  pht_2_56 = _RAND_632[1:0];
  _RAND_633 = {1{`RANDOM}};
  pht_2_57 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  pht_2_58 = _RAND_634[1:0];
  _RAND_635 = {1{`RANDOM}};
  pht_2_59 = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  pht_2_60 = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  pht_2_61 = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  pht_2_62 = _RAND_638[1:0];
  _RAND_639 = {1{`RANDOM}};
  pht_2_63 = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  pht_2_64 = _RAND_640[1:0];
  _RAND_641 = {1{`RANDOM}};
  pht_2_65 = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  pht_2_66 = _RAND_642[1:0];
  _RAND_643 = {1{`RANDOM}};
  pht_2_67 = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  pht_2_68 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  pht_2_69 = _RAND_645[1:0];
  _RAND_646 = {1{`RANDOM}};
  pht_2_70 = _RAND_646[1:0];
  _RAND_647 = {1{`RANDOM}};
  pht_2_71 = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  pht_2_72 = _RAND_648[1:0];
  _RAND_649 = {1{`RANDOM}};
  pht_2_73 = _RAND_649[1:0];
  _RAND_650 = {1{`RANDOM}};
  pht_2_74 = _RAND_650[1:0];
  _RAND_651 = {1{`RANDOM}};
  pht_2_75 = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  pht_2_76 = _RAND_652[1:0];
  _RAND_653 = {1{`RANDOM}};
  pht_2_77 = _RAND_653[1:0];
  _RAND_654 = {1{`RANDOM}};
  pht_2_78 = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  pht_2_79 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  pht_2_80 = _RAND_656[1:0];
  _RAND_657 = {1{`RANDOM}};
  pht_2_81 = _RAND_657[1:0];
  _RAND_658 = {1{`RANDOM}};
  pht_2_82 = _RAND_658[1:0];
  _RAND_659 = {1{`RANDOM}};
  pht_2_83 = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  pht_2_84 = _RAND_660[1:0];
  _RAND_661 = {1{`RANDOM}};
  pht_2_85 = _RAND_661[1:0];
  _RAND_662 = {1{`RANDOM}};
  pht_2_86 = _RAND_662[1:0];
  _RAND_663 = {1{`RANDOM}};
  pht_2_87 = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  pht_2_88 = _RAND_664[1:0];
  _RAND_665 = {1{`RANDOM}};
  pht_2_89 = _RAND_665[1:0];
  _RAND_666 = {1{`RANDOM}};
  pht_2_90 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  pht_2_91 = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  pht_2_92 = _RAND_668[1:0];
  _RAND_669 = {1{`RANDOM}};
  pht_2_93 = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  pht_2_94 = _RAND_670[1:0];
  _RAND_671 = {1{`RANDOM}};
  pht_2_95 = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  pht_2_96 = _RAND_672[1:0];
  _RAND_673 = {1{`RANDOM}};
  pht_2_97 = _RAND_673[1:0];
  _RAND_674 = {1{`RANDOM}};
  pht_2_98 = _RAND_674[1:0];
  _RAND_675 = {1{`RANDOM}};
  pht_2_99 = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  pht_2_100 = _RAND_676[1:0];
  _RAND_677 = {1{`RANDOM}};
  pht_2_101 = _RAND_677[1:0];
  _RAND_678 = {1{`RANDOM}};
  pht_2_102 = _RAND_678[1:0];
  _RAND_679 = {1{`RANDOM}};
  pht_2_103 = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  pht_2_104 = _RAND_680[1:0];
  _RAND_681 = {1{`RANDOM}};
  pht_2_105 = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  pht_2_106 = _RAND_682[1:0];
  _RAND_683 = {1{`RANDOM}};
  pht_2_107 = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  pht_2_108 = _RAND_684[1:0];
  _RAND_685 = {1{`RANDOM}};
  pht_2_109 = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  pht_2_110 = _RAND_686[1:0];
  _RAND_687 = {1{`RANDOM}};
  pht_2_111 = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  pht_2_112 = _RAND_688[1:0];
  _RAND_689 = {1{`RANDOM}};
  pht_2_113 = _RAND_689[1:0];
  _RAND_690 = {1{`RANDOM}};
  pht_2_114 = _RAND_690[1:0];
  _RAND_691 = {1{`RANDOM}};
  pht_2_115 = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  pht_2_116 = _RAND_692[1:0];
  _RAND_693 = {1{`RANDOM}};
  pht_2_117 = _RAND_693[1:0];
  _RAND_694 = {1{`RANDOM}};
  pht_2_118 = _RAND_694[1:0];
  _RAND_695 = {1{`RANDOM}};
  pht_2_119 = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  pht_2_120 = _RAND_696[1:0];
  _RAND_697 = {1{`RANDOM}};
  pht_2_121 = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  pht_2_122 = _RAND_698[1:0];
  _RAND_699 = {1{`RANDOM}};
  pht_2_123 = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  pht_2_124 = _RAND_700[1:0];
  _RAND_701 = {1{`RANDOM}};
  pht_2_125 = _RAND_701[1:0];
  _RAND_702 = {1{`RANDOM}};
  pht_2_126 = _RAND_702[1:0];
  _RAND_703 = {1{`RANDOM}};
  pht_2_127 = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  pht_2_128 = _RAND_704[1:0];
  _RAND_705 = {1{`RANDOM}};
  pht_2_129 = _RAND_705[1:0];
  _RAND_706 = {1{`RANDOM}};
  pht_2_130 = _RAND_706[1:0];
  _RAND_707 = {1{`RANDOM}};
  pht_2_131 = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  pht_2_132 = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  pht_2_133 = _RAND_709[1:0];
  _RAND_710 = {1{`RANDOM}};
  pht_2_134 = _RAND_710[1:0];
  _RAND_711 = {1{`RANDOM}};
  pht_2_135 = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  pht_2_136 = _RAND_712[1:0];
  _RAND_713 = {1{`RANDOM}};
  pht_2_137 = _RAND_713[1:0];
  _RAND_714 = {1{`RANDOM}};
  pht_2_138 = _RAND_714[1:0];
  _RAND_715 = {1{`RANDOM}};
  pht_2_139 = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  pht_2_140 = _RAND_716[1:0];
  _RAND_717 = {1{`RANDOM}};
  pht_2_141 = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  pht_2_142 = _RAND_718[1:0];
  _RAND_719 = {1{`RANDOM}};
  pht_2_143 = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  pht_2_144 = _RAND_720[1:0];
  _RAND_721 = {1{`RANDOM}};
  pht_2_145 = _RAND_721[1:0];
  _RAND_722 = {1{`RANDOM}};
  pht_2_146 = _RAND_722[1:0];
  _RAND_723 = {1{`RANDOM}};
  pht_2_147 = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  pht_2_148 = _RAND_724[1:0];
  _RAND_725 = {1{`RANDOM}};
  pht_2_149 = _RAND_725[1:0];
  _RAND_726 = {1{`RANDOM}};
  pht_2_150 = _RAND_726[1:0];
  _RAND_727 = {1{`RANDOM}};
  pht_2_151 = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  pht_2_152 = _RAND_728[1:0];
  _RAND_729 = {1{`RANDOM}};
  pht_2_153 = _RAND_729[1:0];
  _RAND_730 = {1{`RANDOM}};
  pht_2_154 = _RAND_730[1:0];
  _RAND_731 = {1{`RANDOM}};
  pht_2_155 = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  pht_2_156 = _RAND_732[1:0];
  _RAND_733 = {1{`RANDOM}};
  pht_2_157 = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  pht_2_158 = _RAND_734[1:0];
  _RAND_735 = {1{`RANDOM}};
  pht_2_159 = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  pht_2_160 = _RAND_736[1:0];
  _RAND_737 = {1{`RANDOM}};
  pht_2_161 = _RAND_737[1:0];
  _RAND_738 = {1{`RANDOM}};
  pht_2_162 = _RAND_738[1:0];
  _RAND_739 = {1{`RANDOM}};
  pht_2_163 = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  pht_2_164 = _RAND_740[1:0];
  _RAND_741 = {1{`RANDOM}};
  pht_2_165 = _RAND_741[1:0];
  _RAND_742 = {1{`RANDOM}};
  pht_2_166 = _RAND_742[1:0];
  _RAND_743 = {1{`RANDOM}};
  pht_2_167 = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  pht_2_168 = _RAND_744[1:0];
  _RAND_745 = {1{`RANDOM}};
  pht_2_169 = _RAND_745[1:0];
  _RAND_746 = {1{`RANDOM}};
  pht_2_170 = _RAND_746[1:0];
  _RAND_747 = {1{`RANDOM}};
  pht_2_171 = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  pht_2_172 = _RAND_748[1:0];
  _RAND_749 = {1{`RANDOM}};
  pht_2_173 = _RAND_749[1:0];
  _RAND_750 = {1{`RANDOM}};
  pht_2_174 = _RAND_750[1:0];
  _RAND_751 = {1{`RANDOM}};
  pht_2_175 = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  pht_2_176 = _RAND_752[1:0];
  _RAND_753 = {1{`RANDOM}};
  pht_2_177 = _RAND_753[1:0];
  _RAND_754 = {1{`RANDOM}};
  pht_2_178 = _RAND_754[1:0];
  _RAND_755 = {1{`RANDOM}};
  pht_2_179 = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  pht_2_180 = _RAND_756[1:0];
  _RAND_757 = {1{`RANDOM}};
  pht_2_181 = _RAND_757[1:0];
  _RAND_758 = {1{`RANDOM}};
  pht_2_182 = _RAND_758[1:0];
  _RAND_759 = {1{`RANDOM}};
  pht_2_183 = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  pht_2_184 = _RAND_760[1:0];
  _RAND_761 = {1{`RANDOM}};
  pht_2_185 = _RAND_761[1:0];
  _RAND_762 = {1{`RANDOM}};
  pht_2_186 = _RAND_762[1:0];
  _RAND_763 = {1{`RANDOM}};
  pht_2_187 = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  pht_2_188 = _RAND_764[1:0];
  _RAND_765 = {1{`RANDOM}};
  pht_2_189 = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  pht_2_190 = _RAND_766[1:0];
  _RAND_767 = {1{`RANDOM}};
  pht_2_191 = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  pht_2_192 = _RAND_768[1:0];
  _RAND_769 = {1{`RANDOM}};
  pht_2_193 = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  pht_2_194 = _RAND_770[1:0];
  _RAND_771 = {1{`RANDOM}};
  pht_2_195 = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  pht_2_196 = _RAND_772[1:0];
  _RAND_773 = {1{`RANDOM}};
  pht_2_197 = _RAND_773[1:0];
  _RAND_774 = {1{`RANDOM}};
  pht_2_198 = _RAND_774[1:0];
  _RAND_775 = {1{`RANDOM}};
  pht_2_199 = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  pht_2_200 = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  pht_2_201 = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  pht_2_202 = _RAND_778[1:0];
  _RAND_779 = {1{`RANDOM}};
  pht_2_203 = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  pht_2_204 = _RAND_780[1:0];
  _RAND_781 = {1{`RANDOM}};
  pht_2_205 = _RAND_781[1:0];
  _RAND_782 = {1{`RANDOM}};
  pht_2_206 = _RAND_782[1:0];
  _RAND_783 = {1{`RANDOM}};
  pht_2_207 = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  pht_2_208 = _RAND_784[1:0];
  _RAND_785 = {1{`RANDOM}};
  pht_2_209 = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  pht_2_210 = _RAND_786[1:0];
  _RAND_787 = {1{`RANDOM}};
  pht_2_211 = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  pht_2_212 = _RAND_788[1:0];
  _RAND_789 = {1{`RANDOM}};
  pht_2_213 = _RAND_789[1:0];
  _RAND_790 = {1{`RANDOM}};
  pht_2_214 = _RAND_790[1:0];
  _RAND_791 = {1{`RANDOM}};
  pht_2_215 = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  pht_2_216 = _RAND_792[1:0];
  _RAND_793 = {1{`RANDOM}};
  pht_2_217 = _RAND_793[1:0];
  _RAND_794 = {1{`RANDOM}};
  pht_2_218 = _RAND_794[1:0];
  _RAND_795 = {1{`RANDOM}};
  pht_2_219 = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  pht_2_220 = _RAND_796[1:0];
  _RAND_797 = {1{`RANDOM}};
  pht_2_221 = _RAND_797[1:0];
  _RAND_798 = {1{`RANDOM}};
  pht_2_222 = _RAND_798[1:0];
  _RAND_799 = {1{`RANDOM}};
  pht_2_223 = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  pht_2_224 = _RAND_800[1:0];
  _RAND_801 = {1{`RANDOM}};
  pht_2_225 = _RAND_801[1:0];
  _RAND_802 = {1{`RANDOM}};
  pht_2_226 = _RAND_802[1:0];
  _RAND_803 = {1{`RANDOM}};
  pht_2_227 = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  pht_2_228 = _RAND_804[1:0];
  _RAND_805 = {1{`RANDOM}};
  pht_2_229 = _RAND_805[1:0];
  _RAND_806 = {1{`RANDOM}};
  pht_2_230 = _RAND_806[1:0];
  _RAND_807 = {1{`RANDOM}};
  pht_2_231 = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  pht_2_232 = _RAND_808[1:0];
  _RAND_809 = {1{`RANDOM}};
  pht_2_233 = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  pht_2_234 = _RAND_810[1:0];
  _RAND_811 = {1{`RANDOM}};
  pht_2_235 = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  pht_2_236 = _RAND_812[1:0];
  _RAND_813 = {1{`RANDOM}};
  pht_2_237 = _RAND_813[1:0];
  _RAND_814 = {1{`RANDOM}};
  pht_2_238 = _RAND_814[1:0];
  _RAND_815 = {1{`RANDOM}};
  pht_2_239 = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  pht_2_240 = _RAND_816[1:0];
  _RAND_817 = {1{`RANDOM}};
  pht_2_241 = _RAND_817[1:0];
  _RAND_818 = {1{`RANDOM}};
  pht_2_242 = _RAND_818[1:0];
  _RAND_819 = {1{`RANDOM}};
  pht_2_243 = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  pht_2_244 = _RAND_820[1:0];
  _RAND_821 = {1{`RANDOM}};
  pht_2_245 = _RAND_821[1:0];
  _RAND_822 = {1{`RANDOM}};
  pht_2_246 = _RAND_822[1:0];
  _RAND_823 = {1{`RANDOM}};
  pht_2_247 = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  pht_2_248 = _RAND_824[1:0];
  _RAND_825 = {1{`RANDOM}};
  pht_2_249 = _RAND_825[1:0];
  _RAND_826 = {1{`RANDOM}};
  pht_2_250 = _RAND_826[1:0];
  _RAND_827 = {1{`RANDOM}};
  pht_2_251 = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  pht_2_252 = _RAND_828[1:0];
  _RAND_829 = {1{`RANDOM}};
  pht_2_253 = _RAND_829[1:0];
  _RAND_830 = {1{`RANDOM}};
  pht_2_254 = _RAND_830[1:0];
  _RAND_831 = {1{`RANDOM}};
  pht_2_255 = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  pht_3_0 = _RAND_832[1:0];
  _RAND_833 = {1{`RANDOM}};
  pht_3_1 = _RAND_833[1:0];
  _RAND_834 = {1{`RANDOM}};
  pht_3_2 = _RAND_834[1:0];
  _RAND_835 = {1{`RANDOM}};
  pht_3_3 = _RAND_835[1:0];
  _RAND_836 = {1{`RANDOM}};
  pht_3_4 = _RAND_836[1:0];
  _RAND_837 = {1{`RANDOM}};
  pht_3_5 = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  pht_3_6 = _RAND_838[1:0];
  _RAND_839 = {1{`RANDOM}};
  pht_3_7 = _RAND_839[1:0];
  _RAND_840 = {1{`RANDOM}};
  pht_3_8 = _RAND_840[1:0];
  _RAND_841 = {1{`RANDOM}};
  pht_3_9 = _RAND_841[1:0];
  _RAND_842 = {1{`RANDOM}};
  pht_3_10 = _RAND_842[1:0];
  _RAND_843 = {1{`RANDOM}};
  pht_3_11 = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  pht_3_12 = _RAND_844[1:0];
  _RAND_845 = {1{`RANDOM}};
  pht_3_13 = _RAND_845[1:0];
  _RAND_846 = {1{`RANDOM}};
  pht_3_14 = _RAND_846[1:0];
  _RAND_847 = {1{`RANDOM}};
  pht_3_15 = _RAND_847[1:0];
  _RAND_848 = {1{`RANDOM}};
  pht_3_16 = _RAND_848[1:0];
  _RAND_849 = {1{`RANDOM}};
  pht_3_17 = _RAND_849[1:0];
  _RAND_850 = {1{`RANDOM}};
  pht_3_18 = _RAND_850[1:0];
  _RAND_851 = {1{`RANDOM}};
  pht_3_19 = _RAND_851[1:0];
  _RAND_852 = {1{`RANDOM}};
  pht_3_20 = _RAND_852[1:0];
  _RAND_853 = {1{`RANDOM}};
  pht_3_21 = _RAND_853[1:0];
  _RAND_854 = {1{`RANDOM}};
  pht_3_22 = _RAND_854[1:0];
  _RAND_855 = {1{`RANDOM}};
  pht_3_23 = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  pht_3_24 = _RAND_856[1:0];
  _RAND_857 = {1{`RANDOM}};
  pht_3_25 = _RAND_857[1:0];
  _RAND_858 = {1{`RANDOM}};
  pht_3_26 = _RAND_858[1:0];
  _RAND_859 = {1{`RANDOM}};
  pht_3_27 = _RAND_859[1:0];
  _RAND_860 = {1{`RANDOM}};
  pht_3_28 = _RAND_860[1:0];
  _RAND_861 = {1{`RANDOM}};
  pht_3_29 = _RAND_861[1:0];
  _RAND_862 = {1{`RANDOM}};
  pht_3_30 = _RAND_862[1:0];
  _RAND_863 = {1{`RANDOM}};
  pht_3_31 = _RAND_863[1:0];
  _RAND_864 = {1{`RANDOM}};
  pht_3_32 = _RAND_864[1:0];
  _RAND_865 = {1{`RANDOM}};
  pht_3_33 = _RAND_865[1:0];
  _RAND_866 = {1{`RANDOM}};
  pht_3_34 = _RAND_866[1:0];
  _RAND_867 = {1{`RANDOM}};
  pht_3_35 = _RAND_867[1:0];
  _RAND_868 = {1{`RANDOM}};
  pht_3_36 = _RAND_868[1:0];
  _RAND_869 = {1{`RANDOM}};
  pht_3_37 = _RAND_869[1:0];
  _RAND_870 = {1{`RANDOM}};
  pht_3_38 = _RAND_870[1:0];
  _RAND_871 = {1{`RANDOM}};
  pht_3_39 = _RAND_871[1:0];
  _RAND_872 = {1{`RANDOM}};
  pht_3_40 = _RAND_872[1:0];
  _RAND_873 = {1{`RANDOM}};
  pht_3_41 = _RAND_873[1:0];
  _RAND_874 = {1{`RANDOM}};
  pht_3_42 = _RAND_874[1:0];
  _RAND_875 = {1{`RANDOM}};
  pht_3_43 = _RAND_875[1:0];
  _RAND_876 = {1{`RANDOM}};
  pht_3_44 = _RAND_876[1:0];
  _RAND_877 = {1{`RANDOM}};
  pht_3_45 = _RAND_877[1:0];
  _RAND_878 = {1{`RANDOM}};
  pht_3_46 = _RAND_878[1:0];
  _RAND_879 = {1{`RANDOM}};
  pht_3_47 = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  pht_3_48 = _RAND_880[1:0];
  _RAND_881 = {1{`RANDOM}};
  pht_3_49 = _RAND_881[1:0];
  _RAND_882 = {1{`RANDOM}};
  pht_3_50 = _RAND_882[1:0];
  _RAND_883 = {1{`RANDOM}};
  pht_3_51 = _RAND_883[1:0];
  _RAND_884 = {1{`RANDOM}};
  pht_3_52 = _RAND_884[1:0];
  _RAND_885 = {1{`RANDOM}};
  pht_3_53 = _RAND_885[1:0];
  _RAND_886 = {1{`RANDOM}};
  pht_3_54 = _RAND_886[1:0];
  _RAND_887 = {1{`RANDOM}};
  pht_3_55 = _RAND_887[1:0];
  _RAND_888 = {1{`RANDOM}};
  pht_3_56 = _RAND_888[1:0];
  _RAND_889 = {1{`RANDOM}};
  pht_3_57 = _RAND_889[1:0];
  _RAND_890 = {1{`RANDOM}};
  pht_3_58 = _RAND_890[1:0];
  _RAND_891 = {1{`RANDOM}};
  pht_3_59 = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  pht_3_60 = _RAND_892[1:0];
  _RAND_893 = {1{`RANDOM}};
  pht_3_61 = _RAND_893[1:0];
  _RAND_894 = {1{`RANDOM}};
  pht_3_62 = _RAND_894[1:0];
  _RAND_895 = {1{`RANDOM}};
  pht_3_63 = _RAND_895[1:0];
  _RAND_896 = {1{`RANDOM}};
  pht_3_64 = _RAND_896[1:0];
  _RAND_897 = {1{`RANDOM}};
  pht_3_65 = _RAND_897[1:0];
  _RAND_898 = {1{`RANDOM}};
  pht_3_66 = _RAND_898[1:0];
  _RAND_899 = {1{`RANDOM}};
  pht_3_67 = _RAND_899[1:0];
  _RAND_900 = {1{`RANDOM}};
  pht_3_68 = _RAND_900[1:0];
  _RAND_901 = {1{`RANDOM}};
  pht_3_69 = _RAND_901[1:0];
  _RAND_902 = {1{`RANDOM}};
  pht_3_70 = _RAND_902[1:0];
  _RAND_903 = {1{`RANDOM}};
  pht_3_71 = _RAND_903[1:0];
  _RAND_904 = {1{`RANDOM}};
  pht_3_72 = _RAND_904[1:0];
  _RAND_905 = {1{`RANDOM}};
  pht_3_73 = _RAND_905[1:0];
  _RAND_906 = {1{`RANDOM}};
  pht_3_74 = _RAND_906[1:0];
  _RAND_907 = {1{`RANDOM}};
  pht_3_75 = _RAND_907[1:0];
  _RAND_908 = {1{`RANDOM}};
  pht_3_76 = _RAND_908[1:0];
  _RAND_909 = {1{`RANDOM}};
  pht_3_77 = _RAND_909[1:0];
  _RAND_910 = {1{`RANDOM}};
  pht_3_78 = _RAND_910[1:0];
  _RAND_911 = {1{`RANDOM}};
  pht_3_79 = _RAND_911[1:0];
  _RAND_912 = {1{`RANDOM}};
  pht_3_80 = _RAND_912[1:0];
  _RAND_913 = {1{`RANDOM}};
  pht_3_81 = _RAND_913[1:0];
  _RAND_914 = {1{`RANDOM}};
  pht_3_82 = _RAND_914[1:0];
  _RAND_915 = {1{`RANDOM}};
  pht_3_83 = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  pht_3_84 = _RAND_916[1:0];
  _RAND_917 = {1{`RANDOM}};
  pht_3_85 = _RAND_917[1:0];
  _RAND_918 = {1{`RANDOM}};
  pht_3_86 = _RAND_918[1:0];
  _RAND_919 = {1{`RANDOM}};
  pht_3_87 = _RAND_919[1:0];
  _RAND_920 = {1{`RANDOM}};
  pht_3_88 = _RAND_920[1:0];
  _RAND_921 = {1{`RANDOM}};
  pht_3_89 = _RAND_921[1:0];
  _RAND_922 = {1{`RANDOM}};
  pht_3_90 = _RAND_922[1:0];
  _RAND_923 = {1{`RANDOM}};
  pht_3_91 = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  pht_3_92 = _RAND_924[1:0];
  _RAND_925 = {1{`RANDOM}};
  pht_3_93 = _RAND_925[1:0];
  _RAND_926 = {1{`RANDOM}};
  pht_3_94 = _RAND_926[1:0];
  _RAND_927 = {1{`RANDOM}};
  pht_3_95 = _RAND_927[1:0];
  _RAND_928 = {1{`RANDOM}};
  pht_3_96 = _RAND_928[1:0];
  _RAND_929 = {1{`RANDOM}};
  pht_3_97 = _RAND_929[1:0];
  _RAND_930 = {1{`RANDOM}};
  pht_3_98 = _RAND_930[1:0];
  _RAND_931 = {1{`RANDOM}};
  pht_3_99 = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  pht_3_100 = _RAND_932[1:0];
  _RAND_933 = {1{`RANDOM}};
  pht_3_101 = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  pht_3_102 = _RAND_934[1:0];
  _RAND_935 = {1{`RANDOM}};
  pht_3_103 = _RAND_935[1:0];
  _RAND_936 = {1{`RANDOM}};
  pht_3_104 = _RAND_936[1:0];
  _RAND_937 = {1{`RANDOM}};
  pht_3_105 = _RAND_937[1:0];
  _RAND_938 = {1{`RANDOM}};
  pht_3_106 = _RAND_938[1:0];
  _RAND_939 = {1{`RANDOM}};
  pht_3_107 = _RAND_939[1:0];
  _RAND_940 = {1{`RANDOM}};
  pht_3_108 = _RAND_940[1:0];
  _RAND_941 = {1{`RANDOM}};
  pht_3_109 = _RAND_941[1:0];
  _RAND_942 = {1{`RANDOM}};
  pht_3_110 = _RAND_942[1:0];
  _RAND_943 = {1{`RANDOM}};
  pht_3_111 = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  pht_3_112 = _RAND_944[1:0];
  _RAND_945 = {1{`RANDOM}};
  pht_3_113 = _RAND_945[1:0];
  _RAND_946 = {1{`RANDOM}};
  pht_3_114 = _RAND_946[1:0];
  _RAND_947 = {1{`RANDOM}};
  pht_3_115 = _RAND_947[1:0];
  _RAND_948 = {1{`RANDOM}};
  pht_3_116 = _RAND_948[1:0];
  _RAND_949 = {1{`RANDOM}};
  pht_3_117 = _RAND_949[1:0];
  _RAND_950 = {1{`RANDOM}};
  pht_3_118 = _RAND_950[1:0];
  _RAND_951 = {1{`RANDOM}};
  pht_3_119 = _RAND_951[1:0];
  _RAND_952 = {1{`RANDOM}};
  pht_3_120 = _RAND_952[1:0];
  _RAND_953 = {1{`RANDOM}};
  pht_3_121 = _RAND_953[1:0];
  _RAND_954 = {1{`RANDOM}};
  pht_3_122 = _RAND_954[1:0];
  _RAND_955 = {1{`RANDOM}};
  pht_3_123 = _RAND_955[1:0];
  _RAND_956 = {1{`RANDOM}};
  pht_3_124 = _RAND_956[1:0];
  _RAND_957 = {1{`RANDOM}};
  pht_3_125 = _RAND_957[1:0];
  _RAND_958 = {1{`RANDOM}};
  pht_3_126 = _RAND_958[1:0];
  _RAND_959 = {1{`RANDOM}};
  pht_3_127 = _RAND_959[1:0];
  _RAND_960 = {1{`RANDOM}};
  pht_3_128 = _RAND_960[1:0];
  _RAND_961 = {1{`RANDOM}};
  pht_3_129 = _RAND_961[1:0];
  _RAND_962 = {1{`RANDOM}};
  pht_3_130 = _RAND_962[1:0];
  _RAND_963 = {1{`RANDOM}};
  pht_3_131 = _RAND_963[1:0];
  _RAND_964 = {1{`RANDOM}};
  pht_3_132 = _RAND_964[1:0];
  _RAND_965 = {1{`RANDOM}};
  pht_3_133 = _RAND_965[1:0];
  _RAND_966 = {1{`RANDOM}};
  pht_3_134 = _RAND_966[1:0];
  _RAND_967 = {1{`RANDOM}};
  pht_3_135 = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  pht_3_136 = _RAND_968[1:0];
  _RAND_969 = {1{`RANDOM}};
  pht_3_137 = _RAND_969[1:0];
  _RAND_970 = {1{`RANDOM}};
  pht_3_138 = _RAND_970[1:0];
  _RAND_971 = {1{`RANDOM}};
  pht_3_139 = _RAND_971[1:0];
  _RAND_972 = {1{`RANDOM}};
  pht_3_140 = _RAND_972[1:0];
  _RAND_973 = {1{`RANDOM}};
  pht_3_141 = _RAND_973[1:0];
  _RAND_974 = {1{`RANDOM}};
  pht_3_142 = _RAND_974[1:0];
  _RAND_975 = {1{`RANDOM}};
  pht_3_143 = _RAND_975[1:0];
  _RAND_976 = {1{`RANDOM}};
  pht_3_144 = _RAND_976[1:0];
  _RAND_977 = {1{`RANDOM}};
  pht_3_145 = _RAND_977[1:0];
  _RAND_978 = {1{`RANDOM}};
  pht_3_146 = _RAND_978[1:0];
  _RAND_979 = {1{`RANDOM}};
  pht_3_147 = _RAND_979[1:0];
  _RAND_980 = {1{`RANDOM}};
  pht_3_148 = _RAND_980[1:0];
  _RAND_981 = {1{`RANDOM}};
  pht_3_149 = _RAND_981[1:0];
  _RAND_982 = {1{`RANDOM}};
  pht_3_150 = _RAND_982[1:0];
  _RAND_983 = {1{`RANDOM}};
  pht_3_151 = _RAND_983[1:0];
  _RAND_984 = {1{`RANDOM}};
  pht_3_152 = _RAND_984[1:0];
  _RAND_985 = {1{`RANDOM}};
  pht_3_153 = _RAND_985[1:0];
  _RAND_986 = {1{`RANDOM}};
  pht_3_154 = _RAND_986[1:0];
  _RAND_987 = {1{`RANDOM}};
  pht_3_155 = _RAND_987[1:0];
  _RAND_988 = {1{`RANDOM}};
  pht_3_156 = _RAND_988[1:0];
  _RAND_989 = {1{`RANDOM}};
  pht_3_157 = _RAND_989[1:0];
  _RAND_990 = {1{`RANDOM}};
  pht_3_158 = _RAND_990[1:0];
  _RAND_991 = {1{`RANDOM}};
  pht_3_159 = _RAND_991[1:0];
  _RAND_992 = {1{`RANDOM}};
  pht_3_160 = _RAND_992[1:0];
  _RAND_993 = {1{`RANDOM}};
  pht_3_161 = _RAND_993[1:0];
  _RAND_994 = {1{`RANDOM}};
  pht_3_162 = _RAND_994[1:0];
  _RAND_995 = {1{`RANDOM}};
  pht_3_163 = _RAND_995[1:0];
  _RAND_996 = {1{`RANDOM}};
  pht_3_164 = _RAND_996[1:0];
  _RAND_997 = {1{`RANDOM}};
  pht_3_165 = _RAND_997[1:0];
  _RAND_998 = {1{`RANDOM}};
  pht_3_166 = _RAND_998[1:0];
  _RAND_999 = {1{`RANDOM}};
  pht_3_167 = _RAND_999[1:0];
  _RAND_1000 = {1{`RANDOM}};
  pht_3_168 = _RAND_1000[1:0];
  _RAND_1001 = {1{`RANDOM}};
  pht_3_169 = _RAND_1001[1:0];
  _RAND_1002 = {1{`RANDOM}};
  pht_3_170 = _RAND_1002[1:0];
  _RAND_1003 = {1{`RANDOM}};
  pht_3_171 = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  pht_3_172 = _RAND_1004[1:0];
  _RAND_1005 = {1{`RANDOM}};
  pht_3_173 = _RAND_1005[1:0];
  _RAND_1006 = {1{`RANDOM}};
  pht_3_174 = _RAND_1006[1:0];
  _RAND_1007 = {1{`RANDOM}};
  pht_3_175 = _RAND_1007[1:0];
  _RAND_1008 = {1{`RANDOM}};
  pht_3_176 = _RAND_1008[1:0];
  _RAND_1009 = {1{`RANDOM}};
  pht_3_177 = _RAND_1009[1:0];
  _RAND_1010 = {1{`RANDOM}};
  pht_3_178 = _RAND_1010[1:0];
  _RAND_1011 = {1{`RANDOM}};
  pht_3_179 = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  pht_3_180 = _RAND_1012[1:0];
  _RAND_1013 = {1{`RANDOM}};
  pht_3_181 = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  pht_3_182 = _RAND_1014[1:0];
  _RAND_1015 = {1{`RANDOM}};
  pht_3_183 = _RAND_1015[1:0];
  _RAND_1016 = {1{`RANDOM}};
  pht_3_184 = _RAND_1016[1:0];
  _RAND_1017 = {1{`RANDOM}};
  pht_3_185 = _RAND_1017[1:0];
  _RAND_1018 = {1{`RANDOM}};
  pht_3_186 = _RAND_1018[1:0];
  _RAND_1019 = {1{`RANDOM}};
  pht_3_187 = _RAND_1019[1:0];
  _RAND_1020 = {1{`RANDOM}};
  pht_3_188 = _RAND_1020[1:0];
  _RAND_1021 = {1{`RANDOM}};
  pht_3_189 = _RAND_1021[1:0];
  _RAND_1022 = {1{`RANDOM}};
  pht_3_190 = _RAND_1022[1:0];
  _RAND_1023 = {1{`RANDOM}};
  pht_3_191 = _RAND_1023[1:0];
  _RAND_1024 = {1{`RANDOM}};
  pht_3_192 = _RAND_1024[1:0];
  _RAND_1025 = {1{`RANDOM}};
  pht_3_193 = _RAND_1025[1:0];
  _RAND_1026 = {1{`RANDOM}};
  pht_3_194 = _RAND_1026[1:0];
  _RAND_1027 = {1{`RANDOM}};
  pht_3_195 = _RAND_1027[1:0];
  _RAND_1028 = {1{`RANDOM}};
  pht_3_196 = _RAND_1028[1:0];
  _RAND_1029 = {1{`RANDOM}};
  pht_3_197 = _RAND_1029[1:0];
  _RAND_1030 = {1{`RANDOM}};
  pht_3_198 = _RAND_1030[1:0];
  _RAND_1031 = {1{`RANDOM}};
  pht_3_199 = _RAND_1031[1:0];
  _RAND_1032 = {1{`RANDOM}};
  pht_3_200 = _RAND_1032[1:0];
  _RAND_1033 = {1{`RANDOM}};
  pht_3_201 = _RAND_1033[1:0];
  _RAND_1034 = {1{`RANDOM}};
  pht_3_202 = _RAND_1034[1:0];
  _RAND_1035 = {1{`RANDOM}};
  pht_3_203 = _RAND_1035[1:0];
  _RAND_1036 = {1{`RANDOM}};
  pht_3_204 = _RAND_1036[1:0];
  _RAND_1037 = {1{`RANDOM}};
  pht_3_205 = _RAND_1037[1:0];
  _RAND_1038 = {1{`RANDOM}};
  pht_3_206 = _RAND_1038[1:0];
  _RAND_1039 = {1{`RANDOM}};
  pht_3_207 = _RAND_1039[1:0];
  _RAND_1040 = {1{`RANDOM}};
  pht_3_208 = _RAND_1040[1:0];
  _RAND_1041 = {1{`RANDOM}};
  pht_3_209 = _RAND_1041[1:0];
  _RAND_1042 = {1{`RANDOM}};
  pht_3_210 = _RAND_1042[1:0];
  _RAND_1043 = {1{`RANDOM}};
  pht_3_211 = _RAND_1043[1:0];
  _RAND_1044 = {1{`RANDOM}};
  pht_3_212 = _RAND_1044[1:0];
  _RAND_1045 = {1{`RANDOM}};
  pht_3_213 = _RAND_1045[1:0];
  _RAND_1046 = {1{`RANDOM}};
  pht_3_214 = _RAND_1046[1:0];
  _RAND_1047 = {1{`RANDOM}};
  pht_3_215 = _RAND_1047[1:0];
  _RAND_1048 = {1{`RANDOM}};
  pht_3_216 = _RAND_1048[1:0];
  _RAND_1049 = {1{`RANDOM}};
  pht_3_217 = _RAND_1049[1:0];
  _RAND_1050 = {1{`RANDOM}};
  pht_3_218 = _RAND_1050[1:0];
  _RAND_1051 = {1{`RANDOM}};
  pht_3_219 = _RAND_1051[1:0];
  _RAND_1052 = {1{`RANDOM}};
  pht_3_220 = _RAND_1052[1:0];
  _RAND_1053 = {1{`RANDOM}};
  pht_3_221 = _RAND_1053[1:0];
  _RAND_1054 = {1{`RANDOM}};
  pht_3_222 = _RAND_1054[1:0];
  _RAND_1055 = {1{`RANDOM}};
  pht_3_223 = _RAND_1055[1:0];
  _RAND_1056 = {1{`RANDOM}};
  pht_3_224 = _RAND_1056[1:0];
  _RAND_1057 = {1{`RANDOM}};
  pht_3_225 = _RAND_1057[1:0];
  _RAND_1058 = {1{`RANDOM}};
  pht_3_226 = _RAND_1058[1:0];
  _RAND_1059 = {1{`RANDOM}};
  pht_3_227 = _RAND_1059[1:0];
  _RAND_1060 = {1{`RANDOM}};
  pht_3_228 = _RAND_1060[1:0];
  _RAND_1061 = {1{`RANDOM}};
  pht_3_229 = _RAND_1061[1:0];
  _RAND_1062 = {1{`RANDOM}};
  pht_3_230 = _RAND_1062[1:0];
  _RAND_1063 = {1{`RANDOM}};
  pht_3_231 = _RAND_1063[1:0];
  _RAND_1064 = {1{`RANDOM}};
  pht_3_232 = _RAND_1064[1:0];
  _RAND_1065 = {1{`RANDOM}};
  pht_3_233 = _RAND_1065[1:0];
  _RAND_1066 = {1{`RANDOM}};
  pht_3_234 = _RAND_1066[1:0];
  _RAND_1067 = {1{`RANDOM}};
  pht_3_235 = _RAND_1067[1:0];
  _RAND_1068 = {1{`RANDOM}};
  pht_3_236 = _RAND_1068[1:0];
  _RAND_1069 = {1{`RANDOM}};
  pht_3_237 = _RAND_1069[1:0];
  _RAND_1070 = {1{`RANDOM}};
  pht_3_238 = _RAND_1070[1:0];
  _RAND_1071 = {1{`RANDOM}};
  pht_3_239 = _RAND_1071[1:0];
  _RAND_1072 = {1{`RANDOM}};
  pht_3_240 = _RAND_1072[1:0];
  _RAND_1073 = {1{`RANDOM}};
  pht_3_241 = _RAND_1073[1:0];
  _RAND_1074 = {1{`RANDOM}};
  pht_3_242 = _RAND_1074[1:0];
  _RAND_1075 = {1{`RANDOM}};
  pht_3_243 = _RAND_1075[1:0];
  _RAND_1076 = {1{`RANDOM}};
  pht_3_244 = _RAND_1076[1:0];
  _RAND_1077 = {1{`RANDOM}};
  pht_3_245 = _RAND_1077[1:0];
  _RAND_1078 = {1{`RANDOM}};
  pht_3_246 = _RAND_1078[1:0];
  _RAND_1079 = {1{`RANDOM}};
  pht_3_247 = _RAND_1079[1:0];
  _RAND_1080 = {1{`RANDOM}};
  pht_3_248 = _RAND_1080[1:0];
  _RAND_1081 = {1{`RANDOM}};
  pht_3_249 = _RAND_1081[1:0];
  _RAND_1082 = {1{`RANDOM}};
  pht_3_250 = _RAND_1082[1:0];
  _RAND_1083 = {1{`RANDOM}};
  pht_3_251 = _RAND_1083[1:0];
  _RAND_1084 = {1{`RANDOM}};
  pht_3_252 = _RAND_1084[1:0];
  _RAND_1085 = {1{`RANDOM}};
  pht_3_253 = _RAND_1085[1:0];
  _RAND_1086 = {1{`RANDOM}};
  pht_3_254 = _RAND_1086[1:0];
  _RAND_1087 = {1{`RANDOM}};
  pht_3_255 = _RAND_1087[1:0];
  _RAND_1088 = {1{`RANDOM}};
  pht_4_0 = _RAND_1088[1:0];
  _RAND_1089 = {1{`RANDOM}};
  pht_4_1 = _RAND_1089[1:0];
  _RAND_1090 = {1{`RANDOM}};
  pht_4_2 = _RAND_1090[1:0];
  _RAND_1091 = {1{`RANDOM}};
  pht_4_3 = _RAND_1091[1:0];
  _RAND_1092 = {1{`RANDOM}};
  pht_4_4 = _RAND_1092[1:0];
  _RAND_1093 = {1{`RANDOM}};
  pht_4_5 = _RAND_1093[1:0];
  _RAND_1094 = {1{`RANDOM}};
  pht_4_6 = _RAND_1094[1:0];
  _RAND_1095 = {1{`RANDOM}};
  pht_4_7 = _RAND_1095[1:0];
  _RAND_1096 = {1{`RANDOM}};
  pht_4_8 = _RAND_1096[1:0];
  _RAND_1097 = {1{`RANDOM}};
  pht_4_9 = _RAND_1097[1:0];
  _RAND_1098 = {1{`RANDOM}};
  pht_4_10 = _RAND_1098[1:0];
  _RAND_1099 = {1{`RANDOM}};
  pht_4_11 = _RAND_1099[1:0];
  _RAND_1100 = {1{`RANDOM}};
  pht_4_12 = _RAND_1100[1:0];
  _RAND_1101 = {1{`RANDOM}};
  pht_4_13 = _RAND_1101[1:0];
  _RAND_1102 = {1{`RANDOM}};
  pht_4_14 = _RAND_1102[1:0];
  _RAND_1103 = {1{`RANDOM}};
  pht_4_15 = _RAND_1103[1:0];
  _RAND_1104 = {1{`RANDOM}};
  pht_4_16 = _RAND_1104[1:0];
  _RAND_1105 = {1{`RANDOM}};
  pht_4_17 = _RAND_1105[1:0];
  _RAND_1106 = {1{`RANDOM}};
  pht_4_18 = _RAND_1106[1:0];
  _RAND_1107 = {1{`RANDOM}};
  pht_4_19 = _RAND_1107[1:0];
  _RAND_1108 = {1{`RANDOM}};
  pht_4_20 = _RAND_1108[1:0];
  _RAND_1109 = {1{`RANDOM}};
  pht_4_21 = _RAND_1109[1:0];
  _RAND_1110 = {1{`RANDOM}};
  pht_4_22 = _RAND_1110[1:0];
  _RAND_1111 = {1{`RANDOM}};
  pht_4_23 = _RAND_1111[1:0];
  _RAND_1112 = {1{`RANDOM}};
  pht_4_24 = _RAND_1112[1:0];
  _RAND_1113 = {1{`RANDOM}};
  pht_4_25 = _RAND_1113[1:0];
  _RAND_1114 = {1{`RANDOM}};
  pht_4_26 = _RAND_1114[1:0];
  _RAND_1115 = {1{`RANDOM}};
  pht_4_27 = _RAND_1115[1:0];
  _RAND_1116 = {1{`RANDOM}};
  pht_4_28 = _RAND_1116[1:0];
  _RAND_1117 = {1{`RANDOM}};
  pht_4_29 = _RAND_1117[1:0];
  _RAND_1118 = {1{`RANDOM}};
  pht_4_30 = _RAND_1118[1:0];
  _RAND_1119 = {1{`RANDOM}};
  pht_4_31 = _RAND_1119[1:0];
  _RAND_1120 = {1{`RANDOM}};
  pht_4_32 = _RAND_1120[1:0];
  _RAND_1121 = {1{`RANDOM}};
  pht_4_33 = _RAND_1121[1:0];
  _RAND_1122 = {1{`RANDOM}};
  pht_4_34 = _RAND_1122[1:0];
  _RAND_1123 = {1{`RANDOM}};
  pht_4_35 = _RAND_1123[1:0];
  _RAND_1124 = {1{`RANDOM}};
  pht_4_36 = _RAND_1124[1:0];
  _RAND_1125 = {1{`RANDOM}};
  pht_4_37 = _RAND_1125[1:0];
  _RAND_1126 = {1{`RANDOM}};
  pht_4_38 = _RAND_1126[1:0];
  _RAND_1127 = {1{`RANDOM}};
  pht_4_39 = _RAND_1127[1:0];
  _RAND_1128 = {1{`RANDOM}};
  pht_4_40 = _RAND_1128[1:0];
  _RAND_1129 = {1{`RANDOM}};
  pht_4_41 = _RAND_1129[1:0];
  _RAND_1130 = {1{`RANDOM}};
  pht_4_42 = _RAND_1130[1:0];
  _RAND_1131 = {1{`RANDOM}};
  pht_4_43 = _RAND_1131[1:0];
  _RAND_1132 = {1{`RANDOM}};
  pht_4_44 = _RAND_1132[1:0];
  _RAND_1133 = {1{`RANDOM}};
  pht_4_45 = _RAND_1133[1:0];
  _RAND_1134 = {1{`RANDOM}};
  pht_4_46 = _RAND_1134[1:0];
  _RAND_1135 = {1{`RANDOM}};
  pht_4_47 = _RAND_1135[1:0];
  _RAND_1136 = {1{`RANDOM}};
  pht_4_48 = _RAND_1136[1:0];
  _RAND_1137 = {1{`RANDOM}};
  pht_4_49 = _RAND_1137[1:0];
  _RAND_1138 = {1{`RANDOM}};
  pht_4_50 = _RAND_1138[1:0];
  _RAND_1139 = {1{`RANDOM}};
  pht_4_51 = _RAND_1139[1:0];
  _RAND_1140 = {1{`RANDOM}};
  pht_4_52 = _RAND_1140[1:0];
  _RAND_1141 = {1{`RANDOM}};
  pht_4_53 = _RAND_1141[1:0];
  _RAND_1142 = {1{`RANDOM}};
  pht_4_54 = _RAND_1142[1:0];
  _RAND_1143 = {1{`RANDOM}};
  pht_4_55 = _RAND_1143[1:0];
  _RAND_1144 = {1{`RANDOM}};
  pht_4_56 = _RAND_1144[1:0];
  _RAND_1145 = {1{`RANDOM}};
  pht_4_57 = _RAND_1145[1:0];
  _RAND_1146 = {1{`RANDOM}};
  pht_4_58 = _RAND_1146[1:0];
  _RAND_1147 = {1{`RANDOM}};
  pht_4_59 = _RAND_1147[1:0];
  _RAND_1148 = {1{`RANDOM}};
  pht_4_60 = _RAND_1148[1:0];
  _RAND_1149 = {1{`RANDOM}};
  pht_4_61 = _RAND_1149[1:0];
  _RAND_1150 = {1{`RANDOM}};
  pht_4_62 = _RAND_1150[1:0];
  _RAND_1151 = {1{`RANDOM}};
  pht_4_63 = _RAND_1151[1:0];
  _RAND_1152 = {1{`RANDOM}};
  pht_4_64 = _RAND_1152[1:0];
  _RAND_1153 = {1{`RANDOM}};
  pht_4_65 = _RAND_1153[1:0];
  _RAND_1154 = {1{`RANDOM}};
  pht_4_66 = _RAND_1154[1:0];
  _RAND_1155 = {1{`RANDOM}};
  pht_4_67 = _RAND_1155[1:0];
  _RAND_1156 = {1{`RANDOM}};
  pht_4_68 = _RAND_1156[1:0];
  _RAND_1157 = {1{`RANDOM}};
  pht_4_69 = _RAND_1157[1:0];
  _RAND_1158 = {1{`RANDOM}};
  pht_4_70 = _RAND_1158[1:0];
  _RAND_1159 = {1{`RANDOM}};
  pht_4_71 = _RAND_1159[1:0];
  _RAND_1160 = {1{`RANDOM}};
  pht_4_72 = _RAND_1160[1:0];
  _RAND_1161 = {1{`RANDOM}};
  pht_4_73 = _RAND_1161[1:0];
  _RAND_1162 = {1{`RANDOM}};
  pht_4_74 = _RAND_1162[1:0];
  _RAND_1163 = {1{`RANDOM}};
  pht_4_75 = _RAND_1163[1:0];
  _RAND_1164 = {1{`RANDOM}};
  pht_4_76 = _RAND_1164[1:0];
  _RAND_1165 = {1{`RANDOM}};
  pht_4_77 = _RAND_1165[1:0];
  _RAND_1166 = {1{`RANDOM}};
  pht_4_78 = _RAND_1166[1:0];
  _RAND_1167 = {1{`RANDOM}};
  pht_4_79 = _RAND_1167[1:0];
  _RAND_1168 = {1{`RANDOM}};
  pht_4_80 = _RAND_1168[1:0];
  _RAND_1169 = {1{`RANDOM}};
  pht_4_81 = _RAND_1169[1:0];
  _RAND_1170 = {1{`RANDOM}};
  pht_4_82 = _RAND_1170[1:0];
  _RAND_1171 = {1{`RANDOM}};
  pht_4_83 = _RAND_1171[1:0];
  _RAND_1172 = {1{`RANDOM}};
  pht_4_84 = _RAND_1172[1:0];
  _RAND_1173 = {1{`RANDOM}};
  pht_4_85 = _RAND_1173[1:0];
  _RAND_1174 = {1{`RANDOM}};
  pht_4_86 = _RAND_1174[1:0];
  _RAND_1175 = {1{`RANDOM}};
  pht_4_87 = _RAND_1175[1:0];
  _RAND_1176 = {1{`RANDOM}};
  pht_4_88 = _RAND_1176[1:0];
  _RAND_1177 = {1{`RANDOM}};
  pht_4_89 = _RAND_1177[1:0];
  _RAND_1178 = {1{`RANDOM}};
  pht_4_90 = _RAND_1178[1:0];
  _RAND_1179 = {1{`RANDOM}};
  pht_4_91 = _RAND_1179[1:0];
  _RAND_1180 = {1{`RANDOM}};
  pht_4_92 = _RAND_1180[1:0];
  _RAND_1181 = {1{`RANDOM}};
  pht_4_93 = _RAND_1181[1:0];
  _RAND_1182 = {1{`RANDOM}};
  pht_4_94 = _RAND_1182[1:0];
  _RAND_1183 = {1{`RANDOM}};
  pht_4_95 = _RAND_1183[1:0];
  _RAND_1184 = {1{`RANDOM}};
  pht_4_96 = _RAND_1184[1:0];
  _RAND_1185 = {1{`RANDOM}};
  pht_4_97 = _RAND_1185[1:0];
  _RAND_1186 = {1{`RANDOM}};
  pht_4_98 = _RAND_1186[1:0];
  _RAND_1187 = {1{`RANDOM}};
  pht_4_99 = _RAND_1187[1:0];
  _RAND_1188 = {1{`RANDOM}};
  pht_4_100 = _RAND_1188[1:0];
  _RAND_1189 = {1{`RANDOM}};
  pht_4_101 = _RAND_1189[1:0];
  _RAND_1190 = {1{`RANDOM}};
  pht_4_102 = _RAND_1190[1:0];
  _RAND_1191 = {1{`RANDOM}};
  pht_4_103 = _RAND_1191[1:0];
  _RAND_1192 = {1{`RANDOM}};
  pht_4_104 = _RAND_1192[1:0];
  _RAND_1193 = {1{`RANDOM}};
  pht_4_105 = _RAND_1193[1:0];
  _RAND_1194 = {1{`RANDOM}};
  pht_4_106 = _RAND_1194[1:0];
  _RAND_1195 = {1{`RANDOM}};
  pht_4_107 = _RAND_1195[1:0];
  _RAND_1196 = {1{`RANDOM}};
  pht_4_108 = _RAND_1196[1:0];
  _RAND_1197 = {1{`RANDOM}};
  pht_4_109 = _RAND_1197[1:0];
  _RAND_1198 = {1{`RANDOM}};
  pht_4_110 = _RAND_1198[1:0];
  _RAND_1199 = {1{`RANDOM}};
  pht_4_111 = _RAND_1199[1:0];
  _RAND_1200 = {1{`RANDOM}};
  pht_4_112 = _RAND_1200[1:0];
  _RAND_1201 = {1{`RANDOM}};
  pht_4_113 = _RAND_1201[1:0];
  _RAND_1202 = {1{`RANDOM}};
  pht_4_114 = _RAND_1202[1:0];
  _RAND_1203 = {1{`RANDOM}};
  pht_4_115 = _RAND_1203[1:0];
  _RAND_1204 = {1{`RANDOM}};
  pht_4_116 = _RAND_1204[1:0];
  _RAND_1205 = {1{`RANDOM}};
  pht_4_117 = _RAND_1205[1:0];
  _RAND_1206 = {1{`RANDOM}};
  pht_4_118 = _RAND_1206[1:0];
  _RAND_1207 = {1{`RANDOM}};
  pht_4_119 = _RAND_1207[1:0];
  _RAND_1208 = {1{`RANDOM}};
  pht_4_120 = _RAND_1208[1:0];
  _RAND_1209 = {1{`RANDOM}};
  pht_4_121 = _RAND_1209[1:0];
  _RAND_1210 = {1{`RANDOM}};
  pht_4_122 = _RAND_1210[1:0];
  _RAND_1211 = {1{`RANDOM}};
  pht_4_123 = _RAND_1211[1:0];
  _RAND_1212 = {1{`RANDOM}};
  pht_4_124 = _RAND_1212[1:0];
  _RAND_1213 = {1{`RANDOM}};
  pht_4_125 = _RAND_1213[1:0];
  _RAND_1214 = {1{`RANDOM}};
  pht_4_126 = _RAND_1214[1:0];
  _RAND_1215 = {1{`RANDOM}};
  pht_4_127 = _RAND_1215[1:0];
  _RAND_1216 = {1{`RANDOM}};
  pht_4_128 = _RAND_1216[1:0];
  _RAND_1217 = {1{`RANDOM}};
  pht_4_129 = _RAND_1217[1:0];
  _RAND_1218 = {1{`RANDOM}};
  pht_4_130 = _RAND_1218[1:0];
  _RAND_1219 = {1{`RANDOM}};
  pht_4_131 = _RAND_1219[1:0];
  _RAND_1220 = {1{`RANDOM}};
  pht_4_132 = _RAND_1220[1:0];
  _RAND_1221 = {1{`RANDOM}};
  pht_4_133 = _RAND_1221[1:0];
  _RAND_1222 = {1{`RANDOM}};
  pht_4_134 = _RAND_1222[1:0];
  _RAND_1223 = {1{`RANDOM}};
  pht_4_135 = _RAND_1223[1:0];
  _RAND_1224 = {1{`RANDOM}};
  pht_4_136 = _RAND_1224[1:0];
  _RAND_1225 = {1{`RANDOM}};
  pht_4_137 = _RAND_1225[1:0];
  _RAND_1226 = {1{`RANDOM}};
  pht_4_138 = _RAND_1226[1:0];
  _RAND_1227 = {1{`RANDOM}};
  pht_4_139 = _RAND_1227[1:0];
  _RAND_1228 = {1{`RANDOM}};
  pht_4_140 = _RAND_1228[1:0];
  _RAND_1229 = {1{`RANDOM}};
  pht_4_141 = _RAND_1229[1:0];
  _RAND_1230 = {1{`RANDOM}};
  pht_4_142 = _RAND_1230[1:0];
  _RAND_1231 = {1{`RANDOM}};
  pht_4_143 = _RAND_1231[1:0];
  _RAND_1232 = {1{`RANDOM}};
  pht_4_144 = _RAND_1232[1:0];
  _RAND_1233 = {1{`RANDOM}};
  pht_4_145 = _RAND_1233[1:0];
  _RAND_1234 = {1{`RANDOM}};
  pht_4_146 = _RAND_1234[1:0];
  _RAND_1235 = {1{`RANDOM}};
  pht_4_147 = _RAND_1235[1:0];
  _RAND_1236 = {1{`RANDOM}};
  pht_4_148 = _RAND_1236[1:0];
  _RAND_1237 = {1{`RANDOM}};
  pht_4_149 = _RAND_1237[1:0];
  _RAND_1238 = {1{`RANDOM}};
  pht_4_150 = _RAND_1238[1:0];
  _RAND_1239 = {1{`RANDOM}};
  pht_4_151 = _RAND_1239[1:0];
  _RAND_1240 = {1{`RANDOM}};
  pht_4_152 = _RAND_1240[1:0];
  _RAND_1241 = {1{`RANDOM}};
  pht_4_153 = _RAND_1241[1:0];
  _RAND_1242 = {1{`RANDOM}};
  pht_4_154 = _RAND_1242[1:0];
  _RAND_1243 = {1{`RANDOM}};
  pht_4_155 = _RAND_1243[1:0];
  _RAND_1244 = {1{`RANDOM}};
  pht_4_156 = _RAND_1244[1:0];
  _RAND_1245 = {1{`RANDOM}};
  pht_4_157 = _RAND_1245[1:0];
  _RAND_1246 = {1{`RANDOM}};
  pht_4_158 = _RAND_1246[1:0];
  _RAND_1247 = {1{`RANDOM}};
  pht_4_159 = _RAND_1247[1:0];
  _RAND_1248 = {1{`RANDOM}};
  pht_4_160 = _RAND_1248[1:0];
  _RAND_1249 = {1{`RANDOM}};
  pht_4_161 = _RAND_1249[1:0];
  _RAND_1250 = {1{`RANDOM}};
  pht_4_162 = _RAND_1250[1:0];
  _RAND_1251 = {1{`RANDOM}};
  pht_4_163 = _RAND_1251[1:0];
  _RAND_1252 = {1{`RANDOM}};
  pht_4_164 = _RAND_1252[1:0];
  _RAND_1253 = {1{`RANDOM}};
  pht_4_165 = _RAND_1253[1:0];
  _RAND_1254 = {1{`RANDOM}};
  pht_4_166 = _RAND_1254[1:0];
  _RAND_1255 = {1{`RANDOM}};
  pht_4_167 = _RAND_1255[1:0];
  _RAND_1256 = {1{`RANDOM}};
  pht_4_168 = _RAND_1256[1:0];
  _RAND_1257 = {1{`RANDOM}};
  pht_4_169 = _RAND_1257[1:0];
  _RAND_1258 = {1{`RANDOM}};
  pht_4_170 = _RAND_1258[1:0];
  _RAND_1259 = {1{`RANDOM}};
  pht_4_171 = _RAND_1259[1:0];
  _RAND_1260 = {1{`RANDOM}};
  pht_4_172 = _RAND_1260[1:0];
  _RAND_1261 = {1{`RANDOM}};
  pht_4_173 = _RAND_1261[1:0];
  _RAND_1262 = {1{`RANDOM}};
  pht_4_174 = _RAND_1262[1:0];
  _RAND_1263 = {1{`RANDOM}};
  pht_4_175 = _RAND_1263[1:0];
  _RAND_1264 = {1{`RANDOM}};
  pht_4_176 = _RAND_1264[1:0];
  _RAND_1265 = {1{`RANDOM}};
  pht_4_177 = _RAND_1265[1:0];
  _RAND_1266 = {1{`RANDOM}};
  pht_4_178 = _RAND_1266[1:0];
  _RAND_1267 = {1{`RANDOM}};
  pht_4_179 = _RAND_1267[1:0];
  _RAND_1268 = {1{`RANDOM}};
  pht_4_180 = _RAND_1268[1:0];
  _RAND_1269 = {1{`RANDOM}};
  pht_4_181 = _RAND_1269[1:0];
  _RAND_1270 = {1{`RANDOM}};
  pht_4_182 = _RAND_1270[1:0];
  _RAND_1271 = {1{`RANDOM}};
  pht_4_183 = _RAND_1271[1:0];
  _RAND_1272 = {1{`RANDOM}};
  pht_4_184 = _RAND_1272[1:0];
  _RAND_1273 = {1{`RANDOM}};
  pht_4_185 = _RAND_1273[1:0];
  _RAND_1274 = {1{`RANDOM}};
  pht_4_186 = _RAND_1274[1:0];
  _RAND_1275 = {1{`RANDOM}};
  pht_4_187 = _RAND_1275[1:0];
  _RAND_1276 = {1{`RANDOM}};
  pht_4_188 = _RAND_1276[1:0];
  _RAND_1277 = {1{`RANDOM}};
  pht_4_189 = _RAND_1277[1:0];
  _RAND_1278 = {1{`RANDOM}};
  pht_4_190 = _RAND_1278[1:0];
  _RAND_1279 = {1{`RANDOM}};
  pht_4_191 = _RAND_1279[1:0];
  _RAND_1280 = {1{`RANDOM}};
  pht_4_192 = _RAND_1280[1:0];
  _RAND_1281 = {1{`RANDOM}};
  pht_4_193 = _RAND_1281[1:0];
  _RAND_1282 = {1{`RANDOM}};
  pht_4_194 = _RAND_1282[1:0];
  _RAND_1283 = {1{`RANDOM}};
  pht_4_195 = _RAND_1283[1:0];
  _RAND_1284 = {1{`RANDOM}};
  pht_4_196 = _RAND_1284[1:0];
  _RAND_1285 = {1{`RANDOM}};
  pht_4_197 = _RAND_1285[1:0];
  _RAND_1286 = {1{`RANDOM}};
  pht_4_198 = _RAND_1286[1:0];
  _RAND_1287 = {1{`RANDOM}};
  pht_4_199 = _RAND_1287[1:0];
  _RAND_1288 = {1{`RANDOM}};
  pht_4_200 = _RAND_1288[1:0];
  _RAND_1289 = {1{`RANDOM}};
  pht_4_201 = _RAND_1289[1:0];
  _RAND_1290 = {1{`RANDOM}};
  pht_4_202 = _RAND_1290[1:0];
  _RAND_1291 = {1{`RANDOM}};
  pht_4_203 = _RAND_1291[1:0];
  _RAND_1292 = {1{`RANDOM}};
  pht_4_204 = _RAND_1292[1:0];
  _RAND_1293 = {1{`RANDOM}};
  pht_4_205 = _RAND_1293[1:0];
  _RAND_1294 = {1{`RANDOM}};
  pht_4_206 = _RAND_1294[1:0];
  _RAND_1295 = {1{`RANDOM}};
  pht_4_207 = _RAND_1295[1:0];
  _RAND_1296 = {1{`RANDOM}};
  pht_4_208 = _RAND_1296[1:0];
  _RAND_1297 = {1{`RANDOM}};
  pht_4_209 = _RAND_1297[1:0];
  _RAND_1298 = {1{`RANDOM}};
  pht_4_210 = _RAND_1298[1:0];
  _RAND_1299 = {1{`RANDOM}};
  pht_4_211 = _RAND_1299[1:0];
  _RAND_1300 = {1{`RANDOM}};
  pht_4_212 = _RAND_1300[1:0];
  _RAND_1301 = {1{`RANDOM}};
  pht_4_213 = _RAND_1301[1:0];
  _RAND_1302 = {1{`RANDOM}};
  pht_4_214 = _RAND_1302[1:0];
  _RAND_1303 = {1{`RANDOM}};
  pht_4_215 = _RAND_1303[1:0];
  _RAND_1304 = {1{`RANDOM}};
  pht_4_216 = _RAND_1304[1:0];
  _RAND_1305 = {1{`RANDOM}};
  pht_4_217 = _RAND_1305[1:0];
  _RAND_1306 = {1{`RANDOM}};
  pht_4_218 = _RAND_1306[1:0];
  _RAND_1307 = {1{`RANDOM}};
  pht_4_219 = _RAND_1307[1:0];
  _RAND_1308 = {1{`RANDOM}};
  pht_4_220 = _RAND_1308[1:0];
  _RAND_1309 = {1{`RANDOM}};
  pht_4_221 = _RAND_1309[1:0];
  _RAND_1310 = {1{`RANDOM}};
  pht_4_222 = _RAND_1310[1:0];
  _RAND_1311 = {1{`RANDOM}};
  pht_4_223 = _RAND_1311[1:0];
  _RAND_1312 = {1{`RANDOM}};
  pht_4_224 = _RAND_1312[1:0];
  _RAND_1313 = {1{`RANDOM}};
  pht_4_225 = _RAND_1313[1:0];
  _RAND_1314 = {1{`RANDOM}};
  pht_4_226 = _RAND_1314[1:0];
  _RAND_1315 = {1{`RANDOM}};
  pht_4_227 = _RAND_1315[1:0];
  _RAND_1316 = {1{`RANDOM}};
  pht_4_228 = _RAND_1316[1:0];
  _RAND_1317 = {1{`RANDOM}};
  pht_4_229 = _RAND_1317[1:0];
  _RAND_1318 = {1{`RANDOM}};
  pht_4_230 = _RAND_1318[1:0];
  _RAND_1319 = {1{`RANDOM}};
  pht_4_231 = _RAND_1319[1:0];
  _RAND_1320 = {1{`RANDOM}};
  pht_4_232 = _RAND_1320[1:0];
  _RAND_1321 = {1{`RANDOM}};
  pht_4_233 = _RAND_1321[1:0];
  _RAND_1322 = {1{`RANDOM}};
  pht_4_234 = _RAND_1322[1:0];
  _RAND_1323 = {1{`RANDOM}};
  pht_4_235 = _RAND_1323[1:0];
  _RAND_1324 = {1{`RANDOM}};
  pht_4_236 = _RAND_1324[1:0];
  _RAND_1325 = {1{`RANDOM}};
  pht_4_237 = _RAND_1325[1:0];
  _RAND_1326 = {1{`RANDOM}};
  pht_4_238 = _RAND_1326[1:0];
  _RAND_1327 = {1{`RANDOM}};
  pht_4_239 = _RAND_1327[1:0];
  _RAND_1328 = {1{`RANDOM}};
  pht_4_240 = _RAND_1328[1:0];
  _RAND_1329 = {1{`RANDOM}};
  pht_4_241 = _RAND_1329[1:0];
  _RAND_1330 = {1{`RANDOM}};
  pht_4_242 = _RAND_1330[1:0];
  _RAND_1331 = {1{`RANDOM}};
  pht_4_243 = _RAND_1331[1:0];
  _RAND_1332 = {1{`RANDOM}};
  pht_4_244 = _RAND_1332[1:0];
  _RAND_1333 = {1{`RANDOM}};
  pht_4_245 = _RAND_1333[1:0];
  _RAND_1334 = {1{`RANDOM}};
  pht_4_246 = _RAND_1334[1:0];
  _RAND_1335 = {1{`RANDOM}};
  pht_4_247 = _RAND_1335[1:0];
  _RAND_1336 = {1{`RANDOM}};
  pht_4_248 = _RAND_1336[1:0];
  _RAND_1337 = {1{`RANDOM}};
  pht_4_249 = _RAND_1337[1:0];
  _RAND_1338 = {1{`RANDOM}};
  pht_4_250 = _RAND_1338[1:0];
  _RAND_1339 = {1{`RANDOM}};
  pht_4_251 = _RAND_1339[1:0];
  _RAND_1340 = {1{`RANDOM}};
  pht_4_252 = _RAND_1340[1:0];
  _RAND_1341 = {1{`RANDOM}};
  pht_4_253 = _RAND_1341[1:0];
  _RAND_1342 = {1{`RANDOM}};
  pht_4_254 = _RAND_1342[1:0];
  _RAND_1343 = {1{`RANDOM}};
  pht_4_255 = _RAND_1343[1:0];
  _RAND_1344 = {1{`RANDOM}};
  pht_5_0 = _RAND_1344[1:0];
  _RAND_1345 = {1{`RANDOM}};
  pht_5_1 = _RAND_1345[1:0];
  _RAND_1346 = {1{`RANDOM}};
  pht_5_2 = _RAND_1346[1:0];
  _RAND_1347 = {1{`RANDOM}};
  pht_5_3 = _RAND_1347[1:0];
  _RAND_1348 = {1{`RANDOM}};
  pht_5_4 = _RAND_1348[1:0];
  _RAND_1349 = {1{`RANDOM}};
  pht_5_5 = _RAND_1349[1:0];
  _RAND_1350 = {1{`RANDOM}};
  pht_5_6 = _RAND_1350[1:0];
  _RAND_1351 = {1{`RANDOM}};
  pht_5_7 = _RAND_1351[1:0];
  _RAND_1352 = {1{`RANDOM}};
  pht_5_8 = _RAND_1352[1:0];
  _RAND_1353 = {1{`RANDOM}};
  pht_5_9 = _RAND_1353[1:0];
  _RAND_1354 = {1{`RANDOM}};
  pht_5_10 = _RAND_1354[1:0];
  _RAND_1355 = {1{`RANDOM}};
  pht_5_11 = _RAND_1355[1:0];
  _RAND_1356 = {1{`RANDOM}};
  pht_5_12 = _RAND_1356[1:0];
  _RAND_1357 = {1{`RANDOM}};
  pht_5_13 = _RAND_1357[1:0];
  _RAND_1358 = {1{`RANDOM}};
  pht_5_14 = _RAND_1358[1:0];
  _RAND_1359 = {1{`RANDOM}};
  pht_5_15 = _RAND_1359[1:0];
  _RAND_1360 = {1{`RANDOM}};
  pht_5_16 = _RAND_1360[1:0];
  _RAND_1361 = {1{`RANDOM}};
  pht_5_17 = _RAND_1361[1:0];
  _RAND_1362 = {1{`RANDOM}};
  pht_5_18 = _RAND_1362[1:0];
  _RAND_1363 = {1{`RANDOM}};
  pht_5_19 = _RAND_1363[1:0];
  _RAND_1364 = {1{`RANDOM}};
  pht_5_20 = _RAND_1364[1:0];
  _RAND_1365 = {1{`RANDOM}};
  pht_5_21 = _RAND_1365[1:0];
  _RAND_1366 = {1{`RANDOM}};
  pht_5_22 = _RAND_1366[1:0];
  _RAND_1367 = {1{`RANDOM}};
  pht_5_23 = _RAND_1367[1:0];
  _RAND_1368 = {1{`RANDOM}};
  pht_5_24 = _RAND_1368[1:0];
  _RAND_1369 = {1{`RANDOM}};
  pht_5_25 = _RAND_1369[1:0];
  _RAND_1370 = {1{`RANDOM}};
  pht_5_26 = _RAND_1370[1:0];
  _RAND_1371 = {1{`RANDOM}};
  pht_5_27 = _RAND_1371[1:0];
  _RAND_1372 = {1{`RANDOM}};
  pht_5_28 = _RAND_1372[1:0];
  _RAND_1373 = {1{`RANDOM}};
  pht_5_29 = _RAND_1373[1:0];
  _RAND_1374 = {1{`RANDOM}};
  pht_5_30 = _RAND_1374[1:0];
  _RAND_1375 = {1{`RANDOM}};
  pht_5_31 = _RAND_1375[1:0];
  _RAND_1376 = {1{`RANDOM}};
  pht_5_32 = _RAND_1376[1:0];
  _RAND_1377 = {1{`RANDOM}};
  pht_5_33 = _RAND_1377[1:0];
  _RAND_1378 = {1{`RANDOM}};
  pht_5_34 = _RAND_1378[1:0];
  _RAND_1379 = {1{`RANDOM}};
  pht_5_35 = _RAND_1379[1:0];
  _RAND_1380 = {1{`RANDOM}};
  pht_5_36 = _RAND_1380[1:0];
  _RAND_1381 = {1{`RANDOM}};
  pht_5_37 = _RAND_1381[1:0];
  _RAND_1382 = {1{`RANDOM}};
  pht_5_38 = _RAND_1382[1:0];
  _RAND_1383 = {1{`RANDOM}};
  pht_5_39 = _RAND_1383[1:0];
  _RAND_1384 = {1{`RANDOM}};
  pht_5_40 = _RAND_1384[1:0];
  _RAND_1385 = {1{`RANDOM}};
  pht_5_41 = _RAND_1385[1:0];
  _RAND_1386 = {1{`RANDOM}};
  pht_5_42 = _RAND_1386[1:0];
  _RAND_1387 = {1{`RANDOM}};
  pht_5_43 = _RAND_1387[1:0];
  _RAND_1388 = {1{`RANDOM}};
  pht_5_44 = _RAND_1388[1:0];
  _RAND_1389 = {1{`RANDOM}};
  pht_5_45 = _RAND_1389[1:0];
  _RAND_1390 = {1{`RANDOM}};
  pht_5_46 = _RAND_1390[1:0];
  _RAND_1391 = {1{`RANDOM}};
  pht_5_47 = _RAND_1391[1:0];
  _RAND_1392 = {1{`RANDOM}};
  pht_5_48 = _RAND_1392[1:0];
  _RAND_1393 = {1{`RANDOM}};
  pht_5_49 = _RAND_1393[1:0];
  _RAND_1394 = {1{`RANDOM}};
  pht_5_50 = _RAND_1394[1:0];
  _RAND_1395 = {1{`RANDOM}};
  pht_5_51 = _RAND_1395[1:0];
  _RAND_1396 = {1{`RANDOM}};
  pht_5_52 = _RAND_1396[1:0];
  _RAND_1397 = {1{`RANDOM}};
  pht_5_53 = _RAND_1397[1:0];
  _RAND_1398 = {1{`RANDOM}};
  pht_5_54 = _RAND_1398[1:0];
  _RAND_1399 = {1{`RANDOM}};
  pht_5_55 = _RAND_1399[1:0];
  _RAND_1400 = {1{`RANDOM}};
  pht_5_56 = _RAND_1400[1:0];
  _RAND_1401 = {1{`RANDOM}};
  pht_5_57 = _RAND_1401[1:0];
  _RAND_1402 = {1{`RANDOM}};
  pht_5_58 = _RAND_1402[1:0];
  _RAND_1403 = {1{`RANDOM}};
  pht_5_59 = _RAND_1403[1:0];
  _RAND_1404 = {1{`RANDOM}};
  pht_5_60 = _RAND_1404[1:0];
  _RAND_1405 = {1{`RANDOM}};
  pht_5_61 = _RAND_1405[1:0];
  _RAND_1406 = {1{`RANDOM}};
  pht_5_62 = _RAND_1406[1:0];
  _RAND_1407 = {1{`RANDOM}};
  pht_5_63 = _RAND_1407[1:0];
  _RAND_1408 = {1{`RANDOM}};
  pht_5_64 = _RAND_1408[1:0];
  _RAND_1409 = {1{`RANDOM}};
  pht_5_65 = _RAND_1409[1:0];
  _RAND_1410 = {1{`RANDOM}};
  pht_5_66 = _RAND_1410[1:0];
  _RAND_1411 = {1{`RANDOM}};
  pht_5_67 = _RAND_1411[1:0];
  _RAND_1412 = {1{`RANDOM}};
  pht_5_68 = _RAND_1412[1:0];
  _RAND_1413 = {1{`RANDOM}};
  pht_5_69 = _RAND_1413[1:0];
  _RAND_1414 = {1{`RANDOM}};
  pht_5_70 = _RAND_1414[1:0];
  _RAND_1415 = {1{`RANDOM}};
  pht_5_71 = _RAND_1415[1:0];
  _RAND_1416 = {1{`RANDOM}};
  pht_5_72 = _RAND_1416[1:0];
  _RAND_1417 = {1{`RANDOM}};
  pht_5_73 = _RAND_1417[1:0];
  _RAND_1418 = {1{`RANDOM}};
  pht_5_74 = _RAND_1418[1:0];
  _RAND_1419 = {1{`RANDOM}};
  pht_5_75 = _RAND_1419[1:0];
  _RAND_1420 = {1{`RANDOM}};
  pht_5_76 = _RAND_1420[1:0];
  _RAND_1421 = {1{`RANDOM}};
  pht_5_77 = _RAND_1421[1:0];
  _RAND_1422 = {1{`RANDOM}};
  pht_5_78 = _RAND_1422[1:0];
  _RAND_1423 = {1{`RANDOM}};
  pht_5_79 = _RAND_1423[1:0];
  _RAND_1424 = {1{`RANDOM}};
  pht_5_80 = _RAND_1424[1:0];
  _RAND_1425 = {1{`RANDOM}};
  pht_5_81 = _RAND_1425[1:0];
  _RAND_1426 = {1{`RANDOM}};
  pht_5_82 = _RAND_1426[1:0];
  _RAND_1427 = {1{`RANDOM}};
  pht_5_83 = _RAND_1427[1:0];
  _RAND_1428 = {1{`RANDOM}};
  pht_5_84 = _RAND_1428[1:0];
  _RAND_1429 = {1{`RANDOM}};
  pht_5_85 = _RAND_1429[1:0];
  _RAND_1430 = {1{`RANDOM}};
  pht_5_86 = _RAND_1430[1:0];
  _RAND_1431 = {1{`RANDOM}};
  pht_5_87 = _RAND_1431[1:0];
  _RAND_1432 = {1{`RANDOM}};
  pht_5_88 = _RAND_1432[1:0];
  _RAND_1433 = {1{`RANDOM}};
  pht_5_89 = _RAND_1433[1:0];
  _RAND_1434 = {1{`RANDOM}};
  pht_5_90 = _RAND_1434[1:0];
  _RAND_1435 = {1{`RANDOM}};
  pht_5_91 = _RAND_1435[1:0];
  _RAND_1436 = {1{`RANDOM}};
  pht_5_92 = _RAND_1436[1:0];
  _RAND_1437 = {1{`RANDOM}};
  pht_5_93 = _RAND_1437[1:0];
  _RAND_1438 = {1{`RANDOM}};
  pht_5_94 = _RAND_1438[1:0];
  _RAND_1439 = {1{`RANDOM}};
  pht_5_95 = _RAND_1439[1:0];
  _RAND_1440 = {1{`RANDOM}};
  pht_5_96 = _RAND_1440[1:0];
  _RAND_1441 = {1{`RANDOM}};
  pht_5_97 = _RAND_1441[1:0];
  _RAND_1442 = {1{`RANDOM}};
  pht_5_98 = _RAND_1442[1:0];
  _RAND_1443 = {1{`RANDOM}};
  pht_5_99 = _RAND_1443[1:0];
  _RAND_1444 = {1{`RANDOM}};
  pht_5_100 = _RAND_1444[1:0];
  _RAND_1445 = {1{`RANDOM}};
  pht_5_101 = _RAND_1445[1:0];
  _RAND_1446 = {1{`RANDOM}};
  pht_5_102 = _RAND_1446[1:0];
  _RAND_1447 = {1{`RANDOM}};
  pht_5_103 = _RAND_1447[1:0];
  _RAND_1448 = {1{`RANDOM}};
  pht_5_104 = _RAND_1448[1:0];
  _RAND_1449 = {1{`RANDOM}};
  pht_5_105 = _RAND_1449[1:0];
  _RAND_1450 = {1{`RANDOM}};
  pht_5_106 = _RAND_1450[1:0];
  _RAND_1451 = {1{`RANDOM}};
  pht_5_107 = _RAND_1451[1:0];
  _RAND_1452 = {1{`RANDOM}};
  pht_5_108 = _RAND_1452[1:0];
  _RAND_1453 = {1{`RANDOM}};
  pht_5_109 = _RAND_1453[1:0];
  _RAND_1454 = {1{`RANDOM}};
  pht_5_110 = _RAND_1454[1:0];
  _RAND_1455 = {1{`RANDOM}};
  pht_5_111 = _RAND_1455[1:0];
  _RAND_1456 = {1{`RANDOM}};
  pht_5_112 = _RAND_1456[1:0];
  _RAND_1457 = {1{`RANDOM}};
  pht_5_113 = _RAND_1457[1:0];
  _RAND_1458 = {1{`RANDOM}};
  pht_5_114 = _RAND_1458[1:0];
  _RAND_1459 = {1{`RANDOM}};
  pht_5_115 = _RAND_1459[1:0];
  _RAND_1460 = {1{`RANDOM}};
  pht_5_116 = _RAND_1460[1:0];
  _RAND_1461 = {1{`RANDOM}};
  pht_5_117 = _RAND_1461[1:0];
  _RAND_1462 = {1{`RANDOM}};
  pht_5_118 = _RAND_1462[1:0];
  _RAND_1463 = {1{`RANDOM}};
  pht_5_119 = _RAND_1463[1:0];
  _RAND_1464 = {1{`RANDOM}};
  pht_5_120 = _RAND_1464[1:0];
  _RAND_1465 = {1{`RANDOM}};
  pht_5_121 = _RAND_1465[1:0];
  _RAND_1466 = {1{`RANDOM}};
  pht_5_122 = _RAND_1466[1:0];
  _RAND_1467 = {1{`RANDOM}};
  pht_5_123 = _RAND_1467[1:0];
  _RAND_1468 = {1{`RANDOM}};
  pht_5_124 = _RAND_1468[1:0];
  _RAND_1469 = {1{`RANDOM}};
  pht_5_125 = _RAND_1469[1:0];
  _RAND_1470 = {1{`RANDOM}};
  pht_5_126 = _RAND_1470[1:0];
  _RAND_1471 = {1{`RANDOM}};
  pht_5_127 = _RAND_1471[1:0];
  _RAND_1472 = {1{`RANDOM}};
  pht_5_128 = _RAND_1472[1:0];
  _RAND_1473 = {1{`RANDOM}};
  pht_5_129 = _RAND_1473[1:0];
  _RAND_1474 = {1{`RANDOM}};
  pht_5_130 = _RAND_1474[1:0];
  _RAND_1475 = {1{`RANDOM}};
  pht_5_131 = _RAND_1475[1:0];
  _RAND_1476 = {1{`RANDOM}};
  pht_5_132 = _RAND_1476[1:0];
  _RAND_1477 = {1{`RANDOM}};
  pht_5_133 = _RAND_1477[1:0];
  _RAND_1478 = {1{`RANDOM}};
  pht_5_134 = _RAND_1478[1:0];
  _RAND_1479 = {1{`RANDOM}};
  pht_5_135 = _RAND_1479[1:0];
  _RAND_1480 = {1{`RANDOM}};
  pht_5_136 = _RAND_1480[1:0];
  _RAND_1481 = {1{`RANDOM}};
  pht_5_137 = _RAND_1481[1:0];
  _RAND_1482 = {1{`RANDOM}};
  pht_5_138 = _RAND_1482[1:0];
  _RAND_1483 = {1{`RANDOM}};
  pht_5_139 = _RAND_1483[1:0];
  _RAND_1484 = {1{`RANDOM}};
  pht_5_140 = _RAND_1484[1:0];
  _RAND_1485 = {1{`RANDOM}};
  pht_5_141 = _RAND_1485[1:0];
  _RAND_1486 = {1{`RANDOM}};
  pht_5_142 = _RAND_1486[1:0];
  _RAND_1487 = {1{`RANDOM}};
  pht_5_143 = _RAND_1487[1:0];
  _RAND_1488 = {1{`RANDOM}};
  pht_5_144 = _RAND_1488[1:0];
  _RAND_1489 = {1{`RANDOM}};
  pht_5_145 = _RAND_1489[1:0];
  _RAND_1490 = {1{`RANDOM}};
  pht_5_146 = _RAND_1490[1:0];
  _RAND_1491 = {1{`RANDOM}};
  pht_5_147 = _RAND_1491[1:0];
  _RAND_1492 = {1{`RANDOM}};
  pht_5_148 = _RAND_1492[1:0];
  _RAND_1493 = {1{`RANDOM}};
  pht_5_149 = _RAND_1493[1:0];
  _RAND_1494 = {1{`RANDOM}};
  pht_5_150 = _RAND_1494[1:0];
  _RAND_1495 = {1{`RANDOM}};
  pht_5_151 = _RAND_1495[1:0];
  _RAND_1496 = {1{`RANDOM}};
  pht_5_152 = _RAND_1496[1:0];
  _RAND_1497 = {1{`RANDOM}};
  pht_5_153 = _RAND_1497[1:0];
  _RAND_1498 = {1{`RANDOM}};
  pht_5_154 = _RAND_1498[1:0];
  _RAND_1499 = {1{`RANDOM}};
  pht_5_155 = _RAND_1499[1:0];
  _RAND_1500 = {1{`RANDOM}};
  pht_5_156 = _RAND_1500[1:0];
  _RAND_1501 = {1{`RANDOM}};
  pht_5_157 = _RAND_1501[1:0];
  _RAND_1502 = {1{`RANDOM}};
  pht_5_158 = _RAND_1502[1:0];
  _RAND_1503 = {1{`RANDOM}};
  pht_5_159 = _RAND_1503[1:0];
  _RAND_1504 = {1{`RANDOM}};
  pht_5_160 = _RAND_1504[1:0];
  _RAND_1505 = {1{`RANDOM}};
  pht_5_161 = _RAND_1505[1:0];
  _RAND_1506 = {1{`RANDOM}};
  pht_5_162 = _RAND_1506[1:0];
  _RAND_1507 = {1{`RANDOM}};
  pht_5_163 = _RAND_1507[1:0];
  _RAND_1508 = {1{`RANDOM}};
  pht_5_164 = _RAND_1508[1:0];
  _RAND_1509 = {1{`RANDOM}};
  pht_5_165 = _RAND_1509[1:0];
  _RAND_1510 = {1{`RANDOM}};
  pht_5_166 = _RAND_1510[1:0];
  _RAND_1511 = {1{`RANDOM}};
  pht_5_167 = _RAND_1511[1:0];
  _RAND_1512 = {1{`RANDOM}};
  pht_5_168 = _RAND_1512[1:0];
  _RAND_1513 = {1{`RANDOM}};
  pht_5_169 = _RAND_1513[1:0];
  _RAND_1514 = {1{`RANDOM}};
  pht_5_170 = _RAND_1514[1:0];
  _RAND_1515 = {1{`RANDOM}};
  pht_5_171 = _RAND_1515[1:0];
  _RAND_1516 = {1{`RANDOM}};
  pht_5_172 = _RAND_1516[1:0];
  _RAND_1517 = {1{`RANDOM}};
  pht_5_173 = _RAND_1517[1:0];
  _RAND_1518 = {1{`RANDOM}};
  pht_5_174 = _RAND_1518[1:0];
  _RAND_1519 = {1{`RANDOM}};
  pht_5_175 = _RAND_1519[1:0];
  _RAND_1520 = {1{`RANDOM}};
  pht_5_176 = _RAND_1520[1:0];
  _RAND_1521 = {1{`RANDOM}};
  pht_5_177 = _RAND_1521[1:0];
  _RAND_1522 = {1{`RANDOM}};
  pht_5_178 = _RAND_1522[1:0];
  _RAND_1523 = {1{`RANDOM}};
  pht_5_179 = _RAND_1523[1:0];
  _RAND_1524 = {1{`RANDOM}};
  pht_5_180 = _RAND_1524[1:0];
  _RAND_1525 = {1{`RANDOM}};
  pht_5_181 = _RAND_1525[1:0];
  _RAND_1526 = {1{`RANDOM}};
  pht_5_182 = _RAND_1526[1:0];
  _RAND_1527 = {1{`RANDOM}};
  pht_5_183 = _RAND_1527[1:0];
  _RAND_1528 = {1{`RANDOM}};
  pht_5_184 = _RAND_1528[1:0];
  _RAND_1529 = {1{`RANDOM}};
  pht_5_185 = _RAND_1529[1:0];
  _RAND_1530 = {1{`RANDOM}};
  pht_5_186 = _RAND_1530[1:0];
  _RAND_1531 = {1{`RANDOM}};
  pht_5_187 = _RAND_1531[1:0];
  _RAND_1532 = {1{`RANDOM}};
  pht_5_188 = _RAND_1532[1:0];
  _RAND_1533 = {1{`RANDOM}};
  pht_5_189 = _RAND_1533[1:0];
  _RAND_1534 = {1{`RANDOM}};
  pht_5_190 = _RAND_1534[1:0];
  _RAND_1535 = {1{`RANDOM}};
  pht_5_191 = _RAND_1535[1:0];
  _RAND_1536 = {1{`RANDOM}};
  pht_5_192 = _RAND_1536[1:0];
  _RAND_1537 = {1{`RANDOM}};
  pht_5_193 = _RAND_1537[1:0];
  _RAND_1538 = {1{`RANDOM}};
  pht_5_194 = _RAND_1538[1:0];
  _RAND_1539 = {1{`RANDOM}};
  pht_5_195 = _RAND_1539[1:0];
  _RAND_1540 = {1{`RANDOM}};
  pht_5_196 = _RAND_1540[1:0];
  _RAND_1541 = {1{`RANDOM}};
  pht_5_197 = _RAND_1541[1:0];
  _RAND_1542 = {1{`RANDOM}};
  pht_5_198 = _RAND_1542[1:0];
  _RAND_1543 = {1{`RANDOM}};
  pht_5_199 = _RAND_1543[1:0];
  _RAND_1544 = {1{`RANDOM}};
  pht_5_200 = _RAND_1544[1:0];
  _RAND_1545 = {1{`RANDOM}};
  pht_5_201 = _RAND_1545[1:0];
  _RAND_1546 = {1{`RANDOM}};
  pht_5_202 = _RAND_1546[1:0];
  _RAND_1547 = {1{`RANDOM}};
  pht_5_203 = _RAND_1547[1:0];
  _RAND_1548 = {1{`RANDOM}};
  pht_5_204 = _RAND_1548[1:0];
  _RAND_1549 = {1{`RANDOM}};
  pht_5_205 = _RAND_1549[1:0];
  _RAND_1550 = {1{`RANDOM}};
  pht_5_206 = _RAND_1550[1:0];
  _RAND_1551 = {1{`RANDOM}};
  pht_5_207 = _RAND_1551[1:0];
  _RAND_1552 = {1{`RANDOM}};
  pht_5_208 = _RAND_1552[1:0];
  _RAND_1553 = {1{`RANDOM}};
  pht_5_209 = _RAND_1553[1:0];
  _RAND_1554 = {1{`RANDOM}};
  pht_5_210 = _RAND_1554[1:0];
  _RAND_1555 = {1{`RANDOM}};
  pht_5_211 = _RAND_1555[1:0];
  _RAND_1556 = {1{`RANDOM}};
  pht_5_212 = _RAND_1556[1:0];
  _RAND_1557 = {1{`RANDOM}};
  pht_5_213 = _RAND_1557[1:0];
  _RAND_1558 = {1{`RANDOM}};
  pht_5_214 = _RAND_1558[1:0];
  _RAND_1559 = {1{`RANDOM}};
  pht_5_215 = _RAND_1559[1:0];
  _RAND_1560 = {1{`RANDOM}};
  pht_5_216 = _RAND_1560[1:0];
  _RAND_1561 = {1{`RANDOM}};
  pht_5_217 = _RAND_1561[1:0];
  _RAND_1562 = {1{`RANDOM}};
  pht_5_218 = _RAND_1562[1:0];
  _RAND_1563 = {1{`RANDOM}};
  pht_5_219 = _RAND_1563[1:0];
  _RAND_1564 = {1{`RANDOM}};
  pht_5_220 = _RAND_1564[1:0];
  _RAND_1565 = {1{`RANDOM}};
  pht_5_221 = _RAND_1565[1:0];
  _RAND_1566 = {1{`RANDOM}};
  pht_5_222 = _RAND_1566[1:0];
  _RAND_1567 = {1{`RANDOM}};
  pht_5_223 = _RAND_1567[1:0];
  _RAND_1568 = {1{`RANDOM}};
  pht_5_224 = _RAND_1568[1:0];
  _RAND_1569 = {1{`RANDOM}};
  pht_5_225 = _RAND_1569[1:0];
  _RAND_1570 = {1{`RANDOM}};
  pht_5_226 = _RAND_1570[1:0];
  _RAND_1571 = {1{`RANDOM}};
  pht_5_227 = _RAND_1571[1:0];
  _RAND_1572 = {1{`RANDOM}};
  pht_5_228 = _RAND_1572[1:0];
  _RAND_1573 = {1{`RANDOM}};
  pht_5_229 = _RAND_1573[1:0];
  _RAND_1574 = {1{`RANDOM}};
  pht_5_230 = _RAND_1574[1:0];
  _RAND_1575 = {1{`RANDOM}};
  pht_5_231 = _RAND_1575[1:0];
  _RAND_1576 = {1{`RANDOM}};
  pht_5_232 = _RAND_1576[1:0];
  _RAND_1577 = {1{`RANDOM}};
  pht_5_233 = _RAND_1577[1:0];
  _RAND_1578 = {1{`RANDOM}};
  pht_5_234 = _RAND_1578[1:0];
  _RAND_1579 = {1{`RANDOM}};
  pht_5_235 = _RAND_1579[1:0];
  _RAND_1580 = {1{`RANDOM}};
  pht_5_236 = _RAND_1580[1:0];
  _RAND_1581 = {1{`RANDOM}};
  pht_5_237 = _RAND_1581[1:0];
  _RAND_1582 = {1{`RANDOM}};
  pht_5_238 = _RAND_1582[1:0];
  _RAND_1583 = {1{`RANDOM}};
  pht_5_239 = _RAND_1583[1:0];
  _RAND_1584 = {1{`RANDOM}};
  pht_5_240 = _RAND_1584[1:0];
  _RAND_1585 = {1{`RANDOM}};
  pht_5_241 = _RAND_1585[1:0];
  _RAND_1586 = {1{`RANDOM}};
  pht_5_242 = _RAND_1586[1:0];
  _RAND_1587 = {1{`RANDOM}};
  pht_5_243 = _RAND_1587[1:0];
  _RAND_1588 = {1{`RANDOM}};
  pht_5_244 = _RAND_1588[1:0];
  _RAND_1589 = {1{`RANDOM}};
  pht_5_245 = _RAND_1589[1:0];
  _RAND_1590 = {1{`RANDOM}};
  pht_5_246 = _RAND_1590[1:0];
  _RAND_1591 = {1{`RANDOM}};
  pht_5_247 = _RAND_1591[1:0];
  _RAND_1592 = {1{`RANDOM}};
  pht_5_248 = _RAND_1592[1:0];
  _RAND_1593 = {1{`RANDOM}};
  pht_5_249 = _RAND_1593[1:0];
  _RAND_1594 = {1{`RANDOM}};
  pht_5_250 = _RAND_1594[1:0];
  _RAND_1595 = {1{`RANDOM}};
  pht_5_251 = _RAND_1595[1:0];
  _RAND_1596 = {1{`RANDOM}};
  pht_5_252 = _RAND_1596[1:0];
  _RAND_1597 = {1{`RANDOM}};
  pht_5_253 = _RAND_1597[1:0];
  _RAND_1598 = {1{`RANDOM}};
  pht_5_254 = _RAND_1598[1:0];
  _RAND_1599 = {1{`RANDOM}};
  pht_5_255 = _RAND_1599[1:0];
  _RAND_1600 = {1{`RANDOM}};
  pht_6_0 = _RAND_1600[1:0];
  _RAND_1601 = {1{`RANDOM}};
  pht_6_1 = _RAND_1601[1:0];
  _RAND_1602 = {1{`RANDOM}};
  pht_6_2 = _RAND_1602[1:0];
  _RAND_1603 = {1{`RANDOM}};
  pht_6_3 = _RAND_1603[1:0];
  _RAND_1604 = {1{`RANDOM}};
  pht_6_4 = _RAND_1604[1:0];
  _RAND_1605 = {1{`RANDOM}};
  pht_6_5 = _RAND_1605[1:0];
  _RAND_1606 = {1{`RANDOM}};
  pht_6_6 = _RAND_1606[1:0];
  _RAND_1607 = {1{`RANDOM}};
  pht_6_7 = _RAND_1607[1:0];
  _RAND_1608 = {1{`RANDOM}};
  pht_6_8 = _RAND_1608[1:0];
  _RAND_1609 = {1{`RANDOM}};
  pht_6_9 = _RAND_1609[1:0];
  _RAND_1610 = {1{`RANDOM}};
  pht_6_10 = _RAND_1610[1:0];
  _RAND_1611 = {1{`RANDOM}};
  pht_6_11 = _RAND_1611[1:0];
  _RAND_1612 = {1{`RANDOM}};
  pht_6_12 = _RAND_1612[1:0];
  _RAND_1613 = {1{`RANDOM}};
  pht_6_13 = _RAND_1613[1:0];
  _RAND_1614 = {1{`RANDOM}};
  pht_6_14 = _RAND_1614[1:0];
  _RAND_1615 = {1{`RANDOM}};
  pht_6_15 = _RAND_1615[1:0];
  _RAND_1616 = {1{`RANDOM}};
  pht_6_16 = _RAND_1616[1:0];
  _RAND_1617 = {1{`RANDOM}};
  pht_6_17 = _RAND_1617[1:0];
  _RAND_1618 = {1{`RANDOM}};
  pht_6_18 = _RAND_1618[1:0];
  _RAND_1619 = {1{`RANDOM}};
  pht_6_19 = _RAND_1619[1:0];
  _RAND_1620 = {1{`RANDOM}};
  pht_6_20 = _RAND_1620[1:0];
  _RAND_1621 = {1{`RANDOM}};
  pht_6_21 = _RAND_1621[1:0];
  _RAND_1622 = {1{`RANDOM}};
  pht_6_22 = _RAND_1622[1:0];
  _RAND_1623 = {1{`RANDOM}};
  pht_6_23 = _RAND_1623[1:0];
  _RAND_1624 = {1{`RANDOM}};
  pht_6_24 = _RAND_1624[1:0];
  _RAND_1625 = {1{`RANDOM}};
  pht_6_25 = _RAND_1625[1:0];
  _RAND_1626 = {1{`RANDOM}};
  pht_6_26 = _RAND_1626[1:0];
  _RAND_1627 = {1{`RANDOM}};
  pht_6_27 = _RAND_1627[1:0];
  _RAND_1628 = {1{`RANDOM}};
  pht_6_28 = _RAND_1628[1:0];
  _RAND_1629 = {1{`RANDOM}};
  pht_6_29 = _RAND_1629[1:0];
  _RAND_1630 = {1{`RANDOM}};
  pht_6_30 = _RAND_1630[1:0];
  _RAND_1631 = {1{`RANDOM}};
  pht_6_31 = _RAND_1631[1:0];
  _RAND_1632 = {1{`RANDOM}};
  pht_6_32 = _RAND_1632[1:0];
  _RAND_1633 = {1{`RANDOM}};
  pht_6_33 = _RAND_1633[1:0];
  _RAND_1634 = {1{`RANDOM}};
  pht_6_34 = _RAND_1634[1:0];
  _RAND_1635 = {1{`RANDOM}};
  pht_6_35 = _RAND_1635[1:0];
  _RAND_1636 = {1{`RANDOM}};
  pht_6_36 = _RAND_1636[1:0];
  _RAND_1637 = {1{`RANDOM}};
  pht_6_37 = _RAND_1637[1:0];
  _RAND_1638 = {1{`RANDOM}};
  pht_6_38 = _RAND_1638[1:0];
  _RAND_1639 = {1{`RANDOM}};
  pht_6_39 = _RAND_1639[1:0];
  _RAND_1640 = {1{`RANDOM}};
  pht_6_40 = _RAND_1640[1:0];
  _RAND_1641 = {1{`RANDOM}};
  pht_6_41 = _RAND_1641[1:0];
  _RAND_1642 = {1{`RANDOM}};
  pht_6_42 = _RAND_1642[1:0];
  _RAND_1643 = {1{`RANDOM}};
  pht_6_43 = _RAND_1643[1:0];
  _RAND_1644 = {1{`RANDOM}};
  pht_6_44 = _RAND_1644[1:0];
  _RAND_1645 = {1{`RANDOM}};
  pht_6_45 = _RAND_1645[1:0];
  _RAND_1646 = {1{`RANDOM}};
  pht_6_46 = _RAND_1646[1:0];
  _RAND_1647 = {1{`RANDOM}};
  pht_6_47 = _RAND_1647[1:0];
  _RAND_1648 = {1{`RANDOM}};
  pht_6_48 = _RAND_1648[1:0];
  _RAND_1649 = {1{`RANDOM}};
  pht_6_49 = _RAND_1649[1:0];
  _RAND_1650 = {1{`RANDOM}};
  pht_6_50 = _RAND_1650[1:0];
  _RAND_1651 = {1{`RANDOM}};
  pht_6_51 = _RAND_1651[1:0];
  _RAND_1652 = {1{`RANDOM}};
  pht_6_52 = _RAND_1652[1:0];
  _RAND_1653 = {1{`RANDOM}};
  pht_6_53 = _RAND_1653[1:0];
  _RAND_1654 = {1{`RANDOM}};
  pht_6_54 = _RAND_1654[1:0];
  _RAND_1655 = {1{`RANDOM}};
  pht_6_55 = _RAND_1655[1:0];
  _RAND_1656 = {1{`RANDOM}};
  pht_6_56 = _RAND_1656[1:0];
  _RAND_1657 = {1{`RANDOM}};
  pht_6_57 = _RAND_1657[1:0];
  _RAND_1658 = {1{`RANDOM}};
  pht_6_58 = _RAND_1658[1:0];
  _RAND_1659 = {1{`RANDOM}};
  pht_6_59 = _RAND_1659[1:0];
  _RAND_1660 = {1{`RANDOM}};
  pht_6_60 = _RAND_1660[1:0];
  _RAND_1661 = {1{`RANDOM}};
  pht_6_61 = _RAND_1661[1:0];
  _RAND_1662 = {1{`RANDOM}};
  pht_6_62 = _RAND_1662[1:0];
  _RAND_1663 = {1{`RANDOM}};
  pht_6_63 = _RAND_1663[1:0];
  _RAND_1664 = {1{`RANDOM}};
  pht_6_64 = _RAND_1664[1:0];
  _RAND_1665 = {1{`RANDOM}};
  pht_6_65 = _RAND_1665[1:0];
  _RAND_1666 = {1{`RANDOM}};
  pht_6_66 = _RAND_1666[1:0];
  _RAND_1667 = {1{`RANDOM}};
  pht_6_67 = _RAND_1667[1:0];
  _RAND_1668 = {1{`RANDOM}};
  pht_6_68 = _RAND_1668[1:0];
  _RAND_1669 = {1{`RANDOM}};
  pht_6_69 = _RAND_1669[1:0];
  _RAND_1670 = {1{`RANDOM}};
  pht_6_70 = _RAND_1670[1:0];
  _RAND_1671 = {1{`RANDOM}};
  pht_6_71 = _RAND_1671[1:0];
  _RAND_1672 = {1{`RANDOM}};
  pht_6_72 = _RAND_1672[1:0];
  _RAND_1673 = {1{`RANDOM}};
  pht_6_73 = _RAND_1673[1:0];
  _RAND_1674 = {1{`RANDOM}};
  pht_6_74 = _RAND_1674[1:0];
  _RAND_1675 = {1{`RANDOM}};
  pht_6_75 = _RAND_1675[1:0];
  _RAND_1676 = {1{`RANDOM}};
  pht_6_76 = _RAND_1676[1:0];
  _RAND_1677 = {1{`RANDOM}};
  pht_6_77 = _RAND_1677[1:0];
  _RAND_1678 = {1{`RANDOM}};
  pht_6_78 = _RAND_1678[1:0];
  _RAND_1679 = {1{`RANDOM}};
  pht_6_79 = _RAND_1679[1:0];
  _RAND_1680 = {1{`RANDOM}};
  pht_6_80 = _RAND_1680[1:0];
  _RAND_1681 = {1{`RANDOM}};
  pht_6_81 = _RAND_1681[1:0];
  _RAND_1682 = {1{`RANDOM}};
  pht_6_82 = _RAND_1682[1:0];
  _RAND_1683 = {1{`RANDOM}};
  pht_6_83 = _RAND_1683[1:0];
  _RAND_1684 = {1{`RANDOM}};
  pht_6_84 = _RAND_1684[1:0];
  _RAND_1685 = {1{`RANDOM}};
  pht_6_85 = _RAND_1685[1:0];
  _RAND_1686 = {1{`RANDOM}};
  pht_6_86 = _RAND_1686[1:0];
  _RAND_1687 = {1{`RANDOM}};
  pht_6_87 = _RAND_1687[1:0];
  _RAND_1688 = {1{`RANDOM}};
  pht_6_88 = _RAND_1688[1:0];
  _RAND_1689 = {1{`RANDOM}};
  pht_6_89 = _RAND_1689[1:0];
  _RAND_1690 = {1{`RANDOM}};
  pht_6_90 = _RAND_1690[1:0];
  _RAND_1691 = {1{`RANDOM}};
  pht_6_91 = _RAND_1691[1:0];
  _RAND_1692 = {1{`RANDOM}};
  pht_6_92 = _RAND_1692[1:0];
  _RAND_1693 = {1{`RANDOM}};
  pht_6_93 = _RAND_1693[1:0];
  _RAND_1694 = {1{`RANDOM}};
  pht_6_94 = _RAND_1694[1:0];
  _RAND_1695 = {1{`RANDOM}};
  pht_6_95 = _RAND_1695[1:0];
  _RAND_1696 = {1{`RANDOM}};
  pht_6_96 = _RAND_1696[1:0];
  _RAND_1697 = {1{`RANDOM}};
  pht_6_97 = _RAND_1697[1:0];
  _RAND_1698 = {1{`RANDOM}};
  pht_6_98 = _RAND_1698[1:0];
  _RAND_1699 = {1{`RANDOM}};
  pht_6_99 = _RAND_1699[1:0];
  _RAND_1700 = {1{`RANDOM}};
  pht_6_100 = _RAND_1700[1:0];
  _RAND_1701 = {1{`RANDOM}};
  pht_6_101 = _RAND_1701[1:0];
  _RAND_1702 = {1{`RANDOM}};
  pht_6_102 = _RAND_1702[1:0];
  _RAND_1703 = {1{`RANDOM}};
  pht_6_103 = _RAND_1703[1:0];
  _RAND_1704 = {1{`RANDOM}};
  pht_6_104 = _RAND_1704[1:0];
  _RAND_1705 = {1{`RANDOM}};
  pht_6_105 = _RAND_1705[1:0];
  _RAND_1706 = {1{`RANDOM}};
  pht_6_106 = _RAND_1706[1:0];
  _RAND_1707 = {1{`RANDOM}};
  pht_6_107 = _RAND_1707[1:0];
  _RAND_1708 = {1{`RANDOM}};
  pht_6_108 = _RAND_1708[1:0];
  _RAND_1709 = {1{`RANDOM}};
  pht_6_109 = _RAND_1709[1:0];
  _RAND_1710 = {1{`RANDOM}};
  pht_6_110 = _RAND_1710[1:0];
  _RAND_1711 = {1{`RANDOM}};
  pht_6_111 = _RAND_1711[1:0];
  _RAND_1712 = {1{`RANDOM}};
  pht_6_112 = _RAND_1712[1:0];
  _RAND_1713 = {1{`RANDOM}};
  pht_6_113 = _RAND_1713[1:0];
  _RAND_1714 = {1{`RANDOM}};
  pht_6_114 = _RAND_1714[1:0];
  _RAND_1715 = {1{`RANDOM}};
  pht_6_115 = _RAND_1715[1:0];
  _RAND_1716 = {1{`RANDOM}};
  pht_6_116 = _RAND_1716[1:0];
  _RAND_1717 = {1{`RANDOM}};
  pht_6_117 = _RAND_1717[1:0];
  _RAND_1718 = {1{`RANDOM}};
  pht_6_118 = _RAND_1718[1:0];
  _RAND_1719 = {1{`RANDOM}};
  pht_6_119 = _RAND_1719[1:0];
  _RAND_1720 = {1{`RANDOM}};
  pht_6_120 = _RAND_1720[1:0];
  _RAND_1721 = {1{`RANDOM}};
  pht_6_121 = _RAND_1721[1:0];
  _RAND_1722 = {1{`RANDOM}};
  pht_6_122 = _RAND_1722[1:0];
  _RAND_1723 = {1{`RANDOM}};
  pht_6_123 = _RAND_1723[1:0];
  _RAND_1724 = {1{`RANDOM}};
  pht_6_124 = _RAND_1724[1:0];
  _RAND_1725 = {1{`RANDOM}};
  pht_6_125 = _RAND_1725[1:0];
  _RAND_1726 = {1{`RANDOM}};
  pht_6_126 = _RAND_1726[1:0];
  _RAND_1727 = {1{`RANDOM}};
  pht_6_127 = _RAND_1727[1:0];
  _RAND_1728 = {1{`RANDOM}};
  pht_6_128 = _RAND_1728[1:0];
  _RAND_1729 = {1{`RANDOM}};
  pht_6_129 = _RAND_1729[1:0];
  _RAND_1730 = {1{`RANDOM}};
  pht_6_130 = _RAND_1730[1:0];
  _RAND_1731 = {1{`RANDOM}};
  pht_6_131 = _RAND_1731[1:0];
  _RAND_1732 = {1{`RANDOM}};
  pht_6_132 = _RAND_1732[1:0];
  _RAND_1733 = {1{`RANDOM}};
  pht_6_133 = _RAND_1733[1:0];
  _RAND_1734 = {1{`RANDOM}};
  pht_6_134 = _RAND_1734[1:0];
  _RAND_1735 = {1{`RANDOM}};
  pht_6_135 = _RAND_1735[1:0];
  _RAND_1736 = {1{`RANDOM}};
  pht_6_136 = _RAND_1736[1:0];
  _RAND_1737 = {1{`RANDOM}};
  pht_6_137 = _RAND_1737[1:0];
  _RAND_1738 = {1{`RANDOM}};
  pht_6_138 = _RAND_1738[1:0];
  _RAND_1739 = {1{`RANDOM}};
  pht_6_139 = _RAND_1739[1:0];
  _RAND_1740 = {1{`RANDOM}};
  pht_6_140 = _RAND_1740[1:0];
  _RAND_1741 = {1{`RANDOM}};
  pht_6_141 = _RAND_1741[1:0];
  _RAND_1742 = {1{`RANDOM}};
  pht_6_142 = _RAND_1742[1:0];
  _RAND_1743 = {1{`RANDOM}};
  pht_6_143 = _RAND_1743[1:0];
  _RAND_1744 = {1{`RANDOM}};
  pht_6_144 = _RAND_1744[1:0];
  _RAND_1745 = {1{`RANDOM}};
  pht_6_145 = _RAND_1745[1:0];
  _RAND_1746 = {1{`RANDOM}};
  pht_6_146 = _RAND_1746[1:0];
  _RAND_1747 = {1{`RANDOM}};
  pht_6_147 = _RAND_1747[1:0];
  _RAND_1748 = {1{`RANDOM}};
  pht_6_148 = _RAND_1748[1:0];
  _RAND_1749 = {1{`RANDOM}};
  pht_6_149 = _RAND_1749[1:0];
  _RAND_1750 = {1{`RANDOM}};
  pht_6_150 = _RAND_1750[1:0];
  _RAND_1751 = {1{`RANDOM}};
  pht_6_151 = _RAND_1751[1:0];
  _RAND_1752 = {1{`RANDOM}};
  pht_6_152 = _RAND_1752[1:0];
  _RAND_1753 = {1{`RANDOM}};
  pht_6_153 = _RAND_1753[1:0];
  _RAND_1754 = {1{`RANDOM}};
  pht_6_154 = _RAND_1754[1:0];
  _RAND_1755 = {1{`RANDOM}};
  pht_6_155 = _RAND_1755[1:0];
  _RAND_1756 = {1{`RANDOM}};
  pht_6_156 = _RAND_1756[1:0];
  _RAND_1757 = {1{`RANDOM}};
  pht_6_157 = _RAND_1757[1:0];
  _RAND_1758 = {1{`RANDOM}};
  pht_6_158 = _RAND_1758[1:0];
  _RAND_1759 = {1{`RANDOM}};
  pht_6_159 = _RAND_1759[1:0];
  _RAND_1760 = {1{`RANDOM}};
  pht_6_160 = _RAND_1760[1:0];
  _RAND_1761 = {1{`RANDOM}};
  pht_6_161 = _RAND_1761[1:0];
  _RAND_1762 = {1{`RANDOM}};
  pht_6_162 = _RAND_1762[1:0];
  _RAND_1763 = {1{`RANDOM}};
  pht_6_163 = _RAND_1763[1:0];
  _RAND_1764 = {1{`RANDOM}};
  pht_6_164 = _RAND_1764[1:0];
  _RAND_1765 = {1{`RANDOM}};
  pht_6_165 = _RAND_1765[1:0];
  _RAND_1766 = {1{`RANDOM}};
  pht_6_166 = _RAND_1766[1:0];
  _RAND_1767 = {1{`RANDOM}};
  pht_6_167 = _RAND_1767[1:0];
  _RAND_1768 = {1{`RANDOM}};
  pht_6_168 = _RAND_1768[1:0];
  _RAND_1769 = {1{`RANDOM}};
  pht_6_169 = _RAND_1769[1:0];
  _RAND_1770 = {1{`RANDOM}};
  pht_6_170 = _RAND_1770[1:0];
  _RAND_1771 = {1{`RANDOM}};
  pht_6_171 = _RAND_1771[1:0];
  _RAND_1772 = {1{`RANDOM}};
  pht_6_172 = _RAND_1772[1:0];
  _RAND_1773 = {1{`RANDOM}};
  pht_6_173 = _RAND_1773[1:0];
  _RAND_1774 = {1{`RANDOM}};
  pht_6_174 = _RAND_1774[1:0];
  _RAND_1775 = {1{`RANDOM}};
  pht_6_175 = _RAND_1775[1:0];
  _RAND_1776 = {1{`RANDOM}};
  pht_6_176 = _RAND_1776[1:0];
  _RAND_1777 = {1{`RANDOM}};
  pht_6_177 = _RAND_1777[1:0];
  _RAND_1778 = {1{`RANDOM}};
  pht_6_178 = _RAND_1778[1:0];
  _RAND_1779 = {1{`RANDOM}};
  pht_6_179 = _RAND_1779[1:0];
  _RAND_1780 = {1{`RANDOM}};
  pht_6_180 = _RAND_1780[1:0];
  _RAND_1781 = {1{`RANDOM}};
  pht_6_181 = _RAND_1781[1:0];
  _RAND_1782 = {1{`RANDOM}};
  pht_6_182 = _RAND_1782[1:0];
  _RAND_1783 = {1{`RANDOM}};
  pht_6_183 = _RAND_1783[1:0];
  _RAND_1784 = {1{`RANDOM}};
  pht_6_184 = _RAND_1784[1:0];
  _RAND_1785 = {1{`RANDOM}};
  pht_6_185 = _RAND_1785[1:0];
  _RAND_1786 = {1{`RANDOM}};
  pht_6_186 = _RAND_1786[1:0];
  _RAND_1787 = {1{`RANDOM}};
  pht_6_187 = _RAND_1787[1:0];
  _RAND_1788 = {1{`RANDOM}};
  pht_6_188 = _RAND_1788[1:0];
  _RAND_1789 = {1{`RANDOM}};
  pht_6_189 = _RAND_1789[1:0];
  _RAND_1790 = {1{`RANDOM}};
  pht_6_190 = _RAND_1790[1:0];
  _RAND_1791 = {1{`RANDOM}};
  pht_6_191 = _RAND_1791[1:0];
  _RAND_1792 = {1{`RANDOM}};
  pht_6_192 = _RAND_1792[1:0];
  _RAND_1793 = {1{`RANDOM}};
  pht_6_193 = _RAND_1793[1:0];
  _RAND_1794 = {1{`RANDOM}};
  pht_6_194 = _RAND_1794[1:0];
  _RAND_1795 = {1{`RANDOM}};
  pht_6_195 = _RAND_1795[1:0];
  _RAND_1796 = {1{`RANDOM}};
  pht_6_196 = _RAND_1796[1:0];
  _RAND_1797 = {1{`RANDOM}};
  pht_6_197 = _RAND_1797[1:0];
  _RAND_1798 = {1{`RANDOM}};
  pht_6_198 = _RAND_1798[1:0];
  _RAND_1799 = {1{`RANDOM}};
  pht_6_199 = _RAND_1799[1:0];
  _RAND_1800 = {1{`RANDOM}};
  pht_6_200 = _RAND_1800[1:0];
  _RAND_1801 = {1{`RANDOM}};
  pht_6_201 = _RAND_1801[1:0];
  _RAND_1802 = {1{`RANDOM}};
  pht_6_202 = _RAND_1802[1:0];
  _RAND_1803 = {1{`RANDOM}};
  pht_6_203 = _RAND_1803[1:0];
  _RAND_1804 = {1{`RANDOM}};
  pht_6_204 = _RAND_1804[1:0];
  _RAND_1805 = {1{`RANDOM}};
  pht_6_205 = _RAND_1805[1:0];
  _RAND_1806 = {1{`RANDOM}};
  pht_6_206 = _RAND_1806[1:0];
  _RAND_1807 = {1{`RANDOM}};
  pht_6_207 = _RAND_1807[1:0];
  _RAND_1808 = {1{`RANDOM}};
  pht_6_208 = _RAND_1808[1:0];
  _RAND_1809 = {1{`RANDOM}};
  pht_6_209 = _RAND_1809[1:0];
  _RAND_1810 = {1{`RANDOM}};
  pht_6_210 = _RAND_1810[1:0];
  _RAND_1811 = {1{`RANDOM}};
  pht_6_211 = _RAND_1811[1:0];
  _RAND_1812 = {1{`RANDOM}};
  pht_6_212 = _RAND_1812[1:0];
  _RAND_1813 = {1{`RANDOM}};
  pht_6_213 = _RAND_1813[1:0];
  _RAND_1814 = {1{`RANDOM}};
  pht_6_214 = _RAND_1814[1:0];
  _RAND_1815 = {1{`RANDOM}};
  pht_6_215 = _RAND_1815[1:0];
  _RAND_1816 = {1{`RANDOM}};
  pht_6_216 = _RAND_1816[1:0];
  _RAND_1817 = {1{`RANDOM}};
  pht_6_217 = _RAND_1817[1:0];
  _RAND_1818 = {1{`RANDOM}};
  pht_6_218 = _RAND_1818[1:0];
  _RAND_1819 = {1{`RANDOM}};
  pht_6_219 = _RAND_1819[1:0];
  _RAND_1820 = {1{`RANDOM}};
  pht_6_220 = _RAND_1820[1:0];
  _RAND_1821 = {1{`RANDOM}};
  pht_6_221 = _RAND_1821[1:0];
  _RAND_1822 = {1{`RANDOM}};
  pht_6_222 = _RAND_1822[1:0];
  _RAND_1823 = {1{`RANDOM}};
  pht_6_223 = _RAND_1823[1:0];
  _RAND_1824 = {1{`RANDOM}};
  pht_6_224 = _RAND_1824[1:0];
  _RAND_1825 = {1{`RANDOM}};
  pht_6_225 = _RAND_1825[1:0];
  _RAND_1826 = {1{`RANDOM}};
  pht_6_226 = _RAND_1826[1:0];
  _RAND_1827 = {1{`RANDOM}};
  pht_6_227 = _RAND_1827[1:0];
  _RAND_1828 = {1{`RANDOM}};
  pht_6_228 = _RAND_1828[1:0];
  _RAND_1829 = {1{`RANDOM}};
  pht_6_229 = _RAND_1829[1:0];
  _RAND_1830 = {1{`RANDOM}};
  pht_6_230 = _RAND_1830[1:0];
  _RAND_1831 = {1{`RANDOM}};
  pht_6_231 = _RAND_1831[1:0];
  _RAND_1832 = {1{`RANDOM}};
  pht_6_232 = _RAND_1832[1:0];
  _RAND_1833 = {1{`RANDOM}};
  pht_6_233 = _RAND_1833[1:0];
  _RAND_1834 = {1{`RANDOM}};
  pht_6_234 = _RAND_1834[1:0];
  _RAND_1835 = {1{`RANDOM}};
  pht_6_235 = _RAND_1835[1:0];
  _RAND_1836 = {1{`RANDOM}};
  pht_6_236 = _RAND_1836[1:0];
  _RAND_1837 = {1{`RANDOM}};
  pht_6_237 = _RAND_1837[1:0];
  _RAND_1838 = {1{`RANDOM}};
  pht_6_238 = _RAND_1838[1:0];
  _RAND_1839 = {1{`RANDOM}};
  pht_6_239 = _RAND_1839[1:0];
  _RAND_1840 = {1{`RANDOM}};
  pht_6_240 = _RAND_1840[1:0];
  _RAND_1841 = {1{`RANDOM}};
  pht_6_241 = _RAND_1841[1:0];
  _RAND_1842 = {1{`RANDOM}};
  pht_6_242 = _RAND_1842[1:0];
  _RAND_1843 = {1{`RANDOM}};
  pht_6_243 = _RAND_1843[1:0];
  _RAND_1844 = {1{`RANDOM}};
  pht_6_244 = _RAND_1844[1:0];
  _RAND_1845 = {1{`RANDOM}};
  pht_6_245 = _RAND_1845[1:0];
  _RAND_1846 = {1{`RANDOM}};
  pht_6_246 = _RAND_1846[1:0];
  _RAND_1847 = {1{`RANDOM}};
  pht_6_247 = _RAND_1847[1:0];
  _RAND_1848 = {1{`RANDOM}};
  pht_6_248 = _RAND_1848[1:0];
  _RAND_1849 = {1{`RANDOM}};
  pht_6_249 = _RAND_1849[1:0];
  _RAND_1850 = {1{`RANDOM}};
  pht_6_250 = _RAND_1850[1:0];
  _RAND_1851 = {1{`RANDOM}};
  pht_6_251 = _RAND_1851[1:0];
  _RAND_1852 = {1{`RANDOM}};
  pht_6_252 = _RAND_1852[1:0];
  _RAND_1853 = {1{`RANDOM}};
  pht_6_253 = _RAND_1853[1:0];
  _RAND_1854 = {1{`RANDOM}};
  pht_6_254 = _RAND_1854[1:0];
  _RAND_1855 = {1{`RANDOM}};
  pht_6_255 = _RAND_1855[1:0];
  _RAND_1856 = {1{`RANDOM}};
  pht_7_0 = _RAND_1856[1:0];
  _RAND_1857 = {1{`RANDOM}};
  pht_7_1 = _RAND_1857[1:0];
  _RAND_1858 = {1{`RANDOM}};
  pht_7_2 = _RAND_1858[1:0];
  _RAND_1859 = {1{`RANDOM}};
  pht_7_3 = _RAND_1859[1:0];
  _RAND_1860 = {1{`RANDOM}};
  pht_7_4 = _RAND_1860[1:0];
  _RAND_1861 = {1{`RANDOM}};
  pht_7_5 = _RAND_1861[1:0];
  _RAND_1862 = {1{`RANDOM}};
  pht_7_6 = _RAND_1862[1:0];
  _RAND_1863 = {1{`RANDOM}};
  pht_7_7 = _RAND_1863[1:0];
  _RAND_1864 = {1{`RANDOM}};
  pht_7_8 = _RAND_1864[1:0];
  _RAND_1865 = {1{`RANDOM}};
  pht_7_9 = _RAND_1865[1:0];
  _RAND_1866 = {1{`RANDOM}};
  pht_7_10 = _RAND_1866[1:0];
  _RAND_1867 = {1{`RANDOM}};
  pht_7_11 = _RAND_1867[1:0];
  _RAND_1868 = {1{`RANDOM}};
  pht_7_12 = _RAND_1868[1:0];
  _RAND_1869 = {1{`RANDOM}};
  pht_7_13 = _RAND_1869[1:0];
  _RAND_1870 = {1{`RANDOM}};
  pht_7_14 = _RAND_1870[1:0];
  _RAND_1871 = {1{`RANDOM}};
  pht_7_15 = _RAND_1871[1:0];
  _RAND_1872 = {1{`RANDOM}};
  pht_7_16 = _RAND_1872[1:0];
  _RAND_1873 = {1{`RANDOM}};
  pht_7_17 = _RAND_1873[1:0];
  _RAND_1874 = {1{`RANDOM}};
  pht_7_18 = _RAND_1874[1:0];
  _RAND_1875 = {1{`RANDOM}};
  pht_7_19 = _RAND_1875[1:0];
  _RAND_1876 = {1{`RANDOM}};
  pht_7_20 = _RAND_1876[1:0];
  _RAND_1877 = {1{`RANDOM}};
  pht_7_21 = _RAND_1877[1:0];
  _RAND_1878 = {1{`RANDOM}};
  pht_7_22 = _RAND_1878[1:0];
  _RAND_1879 = {1{`RANDOM}};
  pht_7_23 = _RAND_1879[1:0];
  _RAND_1880 = {1{`RANDOM}};
  pht_7_24 = _RAND_1880[1:0];
  _RAND_1881 = {1{`RANDOM}};
  pht_7_25 = _RAND_1881[1:0];
  _RAND_1882 = {1{`RANDOM}};
  pht_7_26 = _RAND_1882[1:0];
  _RAND_1883 = {1{`RANDOM}};
  pht_7_27 = _RAND_1883[1:0];
  _RAND_1884 = {1{`RANDOM}};
  pht_7_28 = _RAND_1884[1:0];
  _RAND_1885 = {1{`RANDOM}};
  pht_7_29 = _RAND_1885[1:0];
  _RAND_1886 = {1{`RANDOM}};
  pht_7_30 = _RAND_1886[1:0];
  _RAND_1887 = {1{`RANDOM}};
  pht_7_31 = _RAND_1887[1:0];
  _RAND_1888 = {1{`RANDOM}};
  pht_7_32 = _RAND_1888[1:0];
  _RAND_1889 = {1{`RANDOM}};
  pht_7_33 = _RAND_1889[1:0];
  _RAND_1890 = {1{`RANDOM}};
  pht_7_34 = _RAND_1890[1:0];
  _RAND_1891 = {1{`RANDOM}};
  pht_7_35 = _RAND_1891[1:0];
  _RAND_1892 = {1{`RANDOM}};
  pht_7_36 = _RAND_1892[1:0];
  _RAND_1893 = {1{`RANDOM}};
  pht_7_37 = _RAND_1893[1:0];
  _RAND_1894 = {1{`RANDOM}};
  pht_7_38 = _RAND_1894[1:0];
  _RAND_1895 = {1{`RANDOM}};
  pht_7_39 = _RAND_1895[1:0];
  _RAND_1896 = {1{`RANDOM}};
  pht_7_40 = _RAND_1896[1:0];
  _RAND_1897 = {1{`RANDOM}};
  pht_7_41 = _RAND_1897[1:0];
  _RAND_1898 = {1{`RANDOM}};
  pht_7_42 = _RAND_1898[1:0];
  _RAND_1899 = {1{`RANDOM}};
  pht_7_43 = _RAND_1899[1:0];
  _RAND_1900 = {1{`RANDOM}};
  pht_7_44 = _RAND_1900[1:0];
  _RAND_1901 = {1{`RANDOM}};
  pht_7_45 = _RAND_1901[1:0];
  _RAND_1902 = {1{`RANDOM}};
  pht_7_46 = _RAND_1902[1:0];
  _RAND_1903 = {1{`RANDOM}};
  pht_7_47 = _RAND_1903[1:0];
  _RAND_1904 = {1{`RANDOM}};
  pht_7_48 = _RAND_1904[1:0];
  _RAND_1905 = {1{`RANDOM}};
  pht_7_49 = _RAND_1905[1:0];
  _RAND_1906 = {1{`RANDOM}};
  pht_7_50 = _RAND_1906[1:0];
  _RAND_1907 = {1{`RANDOM}};
  pht_7_51 = _RAND_1907[1:0];
  _RAND_1908 = {1{`RANDOM}};
  pht_7_52 = _RAND_1908[1:0];
  _RAND_1909 = {1{`RANDOM}};
  pht_7_53 = _RAND_1909[1:0];
  _RAND_1910 = {1{`RANDOM}};
  pht_7_54 = _RAND_1910[1:0];
  _RAND_1911 = {1{`RANDOM}};
  pht_7_55 = _RAND_1911[1:0];
  _RAND_1912 = {1{`RANDOM}};
  pht_7_56 = _RAND_1912[1:0];
  _RAND_1913 = {1{`RANDOM}};
  pht_7_57 = _RAND_1913[1:0];
  _RAND_1914 = {1{`RANDOM}};
  pht_7_58 = _RAND_1914[1:0];
  _RAND_1915 = {1{`RANDOM}};
  pht_7_59 = _RAND_1915[1:0];
  _RAND_1916 = {1{`RANDOM}};
  pht_7_60 = _RAND_1916[1:0];
  _RAND_1917 = {1{`RANDOM}};
  pht_7_61 = _RAND_1917[1:0];
  _RAND_1918 = {1{`RANDOM}};
  pht_7_62 = _RAND_1918[1:0];
  _RAND_1919 = {1{`RANDOM}};
  pht_7_63 = _RAND_1919[1:0];
  _RAND_1920 = {1{`RANDOM}};
  pht_7_64 = _RAND_1920[1:0];
  _RAND_1921 = {1{`RANDOM}};
  pht_7_65 = _RAND_1921[1:0];
  _RAND_1922 = {1{`RANDOM}};
  pht_7_66 = _RAND_1922[1:0];
  _RAND_1923 = {1{`RANDOM}};
  pht_7_67 = _RAND_1923[1:0];
  _RAND_1924 = {1{`RANDOM}};
  pht_7_68 = _RAND_1924[1:0];
  _RAND_1925 = {1{`RANDOM}};
  pht_7_69 = _RAND_1925[1:0];
  _RAND_1926 = {1{`RANDOM}};
  pht_7_70 = _RAND_1926[1:0];
  _RAND_1927 = {1{`RANDOM}};
  pht_7_71 = _RAND_1927[1:0];
  _RAND_1928 = {1{`RANDOM}};
  pht_7_72 = _RAND_1928[1:0];
  _RAND_1929 = {1{`RANDOM}};
  pht_7_73 = _RAND_1929[1:0];
  _RAND_1930 = {1{`RANDOM}};
  pht_7_74 = _RAND_1930[1:0];
  _RAND_1931 = {1{`RANDOM}};
  pht_7_75 = _RAND_1931[1:0];
  _RAND_1932 = {1{`RANDOM}};
  pht_7_76 = _RAND_1932[1:0];
  _RAND_1933 = {1{`RANDOM}};
  pht_7_77 = _RAND_1933[1:0];
  _RAND_1934 = {1{`RANDOM}};
  pht_7_78 = _RAND_1934[1:0];
  _RAND_1935 = {1{`RANDOM}};
  pht_7_79 = _RAND_1935[1:0];
  _RAND_1936 = {1{`RANDOM}};
  pht_7_80 = _RAND_1936[1:0];
  _RAND_1937 = {1{`RANDOM}};
  pht_7_81 = _RAND_1937[1:0];
  _RAND_1938 = {1{`RANDOM}};
  pht_7_82 = _RAND_1938[1:0];
  _RAND_1939 = {1{`RANDOM}};
  pht_7_83 = _RAND_1939[1:0];
  _RAND_1940 = {1{`RANDOM}};
  pht_7_84 = _RAND_1940[1:0];
  _RAND_1941 = {1{`RANDOM}};
  pht_7_85 = _RAND_1941[1:0];
  _RAND_1942 = {1{`RANDOM}};
  pht_7_86 = _RAND_1942[1:0];
  _RAND_1943 = {1{`RANDOM}};
  pht_7_87 = _RAND_1943[1:0];
  _RAND_1944 = {1{`RANDOM}};
  pht_7_88 = _RAND_1944[1:0];
  _RAND_1945 = {1{`RANDOM}};
  pht_7_89 = _RAND_1945[1:0];
  _RAND_1946 = {1{`RANDOM}};
  pht_7_90 = _RAND_1946[1:0];
  _RAND_1947 = {1{`RANDOM}};
  pht_7_91 = _RAND_1947[1:0];
  _RAND_1948 = {1{`RANDOM}};
  pht_7_92 = _RAND_1948[1:0];
  _RAND_1949 = {1{`RANDOM}};
  pht_7_93 = _RAND_1949[1:0];
  _RAND_1950 = {1{`RANDOM}};
  pht_7_94 = _RAND_1950[1:0];
  _RAND_1951 = {1{`RANDOM}};
  pht_7_95 = _RAND_1951[1:0];
  _RAND_1952 = {1{`RANDOM}};
  pht_7_96 = _RAND_1952[1:0];
  _RAND_1953 = {1{`RANDOM}};
  pht_7_97 = _RAND_1953[1:0];
  _RAND_1954 = {1{`RANDOM}};
  pht_7_98 = _RAND_1954[1:0];
  _RAND_1955 = {1{`RANDOM}};
  pht_7_99 = _RAND_1955[1:0];
  _RAND_1956 = {1{`RANDOM}};
  pht_7_100 = _RAND_1956[1:0];
  _RAND_1957 = {1{`RANDOM}};
  pht_7_101 = _RAND_1957[1:0];
  _RAND_1958 = {1{`RANDOM}};
  pht_7_102 = _RAND_1958[1:0];
  _RAND_1959 = {1{`RANDOM}};
  pht_7_103 = _RAND_1959[1:0];
  _RAND_1960 = {1{`RANDOM}};
  pht_7_104 = _RAND_1960[1:0];
  _RAND_1961 = {1{`RANDOM}};
  pht_7_105 = _RAND_1961[1:0];
  _RAND_1962 = {1{`RANDOM}};
  pht_7_106 = _RAND_1962[1:0];
  _RAND_1963 = {1{`RANDOM}};
  pht_7_107 = _RAND_1963[1:0];
  _RAND_1964 = {1{`RANDOM}};
  pht_7_108 = _RAND_1964[1:0];
  _RAND_1965 = {1{`RANDOM}};
  pht_7_109 = _RAND_1965[1:0];
  _RAND_1966 = {1{`RANDOM}};
  pht_7_110 = _RAND_1966[1:0];
  _RAND_1967 = {1{`RANDOM}};
  pht_7_111 = _RAND_1967[1:0];
  _RAND_1968 = {1{`RANDOM}};
  pht_7_112 = _RAND_1968[1:0];
  _RAND_1969 = {1{`RANDOM}};
  pht_7_113 = _RAND_1969[1:0];
  _RAND_1970 = {1{`RANDOM}};
  pht_7_114 = _RAND_1970[1:0];
  _RAND_1971 = {1{`RANDOM}};
  pht_7_115 = _RAND_1971[1:0];
  _RAND_1972 = {1{`RANDOM}};
  pht_7_116 = _RAND_1972[1:0];
  _RAND_1973 = {1{`RANDOM}};
  pht_7_117 = _RAND_1973[1:0];
  _RAND_1974 = {1{`RANDOM}};
  pht_7_118 = _RAND_1974[1:0];
  _RAND_1975 = {1{`RANDOM}};
  pht_7_119 = _RAND_1975[1:0];
  _RAND_1976 = {1{`RANDOM}};
  pht_7_120 = _RAND_1976[1:0];
  _RAND_1977 = {1{`RANDOM}};
  pht_7_121 = _RAND_1977[1:0];
  _RAND_1978 = {1{`RANDOM}};
  pht_7_122 = _RAND_1978[1:0];
  _RAND_1979 = {1{`RANDOM}};
  pht_7_123 = _RAND_1979[1:0];
  _RAND_1980 = {1{`RANDOM}};
  pht_7_124 = _RAND_1980[1:0];
  _RAND_1981 = {1{`RANDOM}};
  pht_7_125 = _RAND_1981[1:0];
  _RAND_1982 = {1{`RANDOM}};
  pht_7_126 = _RAND_1982[1:0];
  _RAND_1983 = {1{`RANDOM}};
  pht_7_127 = _RAND_1983[1:0];
  _RAND_1984 = {1{`RANDOM}};
  pht_7_128 = _RAND_1984[1:0];
  _RAND_1985 = {1{`RANDOM}};
  pht_7_129 = _RAND_1985[1:0];
  _RAND_1986 = {1{`RANDOM}};
  pht_7_130 = _RAND_1986[1:0];
  _RAND_1987 = {1{`RANDOM}};
  pht_7_131 = _RAND_1987[1:0];
  _RAND_1988 = {1{`RANDOM}};
  pht_7_132 = _RAND_1988[1:0];
  _RAND_1989 = {1{`RANDOM}};
  pht_7_133 = _RAND_1989[1:0];
  _RAND_1990 = {1{`RANDOM}};
  pht_7_134 = _RAND_1990[1:0];
  _RAND_1991 = {1{`RANDOM}};
  pht_7_135 = _RAND_1991[1:0];
  _RAND_1992 = {1{`RANDOM}};
  pht_7_136 = _RAND_1992[1:0];
  _RAND_1993 = {1{`RANDOM}};
  pht_7_137 = _RAND_1993[1:0];
  _RAND_1994 = {1{`RANDOM}};
  pht_7_138 = _RAND_1994[1:0];
  _RAND_1995 = {1{`RANDOM}};
  pht_7_139 = _RAND_1995[1:0];
  _RAND_1996 = {1{`RANDOM}};
  pht_7_140 = _RAND_1996[1:0];
  _RAND_1997 = {1{`RANDOM}};
  pht_7_141 = _RAND_1997[1:0];
  _RAND_1998 = {1{`RANDOM}};
  pht_7_142 = _RAND_1998[1:0];
  _RAND_1999 = {1{`RANDOM}};
  pht_7_143 = _RAND_1999[1:0];
  _RAND_2000 = {1{`RANDOM}};
  pht_7_144 = _RAND_2000[1:0];
  _RAND_2001 = {1{`RANDOM}};
  pht_7_145 = _RAND_2001[1:0];
  _RAND_2002 = {1{`RANDOM}};
  pht_7_146 = _RAND_2002[1:0];
  _RAND_2003 = {1{`RANDOM}};
  pht_7_147 = _RAND_2003[1:0];
  _RAND_2004 = {1{`RANDOM}};
  pht_7_148 = _RAND_2004[1:0];
  _RAND_2005 = {1{`RANDOM}};
  pht_7_149 = _RAND_2005[1:0];
  _RAND_2006 = {1{`RANDOM}};
  pht_7_150 = _RAND_2006[1:0];
  _RAND_2007 = {1{`RANDOM}};
  pht_7_151 = _RAND_2007[1:0];
  _RAND_2008 = {1{`RANDOM}};
  pht_7_152 = _RAND_2008[1:0];
  _RAND_2009 = {1{`RANDOM}};
  pht_7_153 = _RAND_2009[1:0];
  _RAND_2010 = {1{`RANDOM}};
  pht_7_154 = _RAND_2010[1:0];
  _RAND_2011 = {1{`RANDOM}};
  pht_7_155 = _RAND_2011[1:0];
  _RAND_2012 = {1{`RANDOM}};
  pht_7_156 = _RAND_2012[1:0];
  _RAND_2013 = {1{`RANDOM}};
  pht_7_157 = _RAND_2013[1:0];
  _RAND_2014 = {1{`RANDOM}};
  pht_7_158 = _RAND_2014[1:0];
  _RAND_2015 = {1{`RANDOM}};
  pht_7_159 = _RAND_2015[1:0];
  _RAND_2016 = {1{`RANDOM}};
  pht_7_160 = _RAND_2016[1:0];
  _RAND_2017 = {1{`RANDOM}};
  pht_7_161 = _RAND_2017[1:0];
  _RAND_2018 = {1{`RANDOM}};
  pht_7_162 = _RAND_2018[1:0];
  _RAND_2019 = {1{`RANDOM}};
  pht_7_163 = _RAND_2019[1:0];
  _RAND_2020 = {1{`RANDOM}};
  pht_7_164 = _RAND_2020[1:0];
  _RAND_2021 = {1{`RANDOM}};
  pht_7_165 = _RAND_2021[1:0];
  _RAND_2022 = {1{`RANDOM}};
  pht_7_166 = _RAND_2022[1:0];
  _RAND_2023 = {1{`RANDOM}};
  pht_7_167 = _RAND_2023[1:0];
  _RAND_2024 = {1{`RANDOM}};
  pht_7_168 = _RAND_2024[1:0];
  _RAND_2025 = {1{`RANDOM}};
  pht_7_169 = _RAND_2025[1:0];
  _RAND_2026 = {1{`RANDOM}};
  pht_7_170 = _RAND_2026[1:0];
  _RAND_2027 = {1{`RANDOM}};
  pht_7_171 = _RAND_2027[1:0];
  _RAND_2028 = {1{`RANDOM}};
  pht_7_172 = _RAND_2028[1:0];
  _RAND_2029 = {1{`RANDOM}};
  pht_7_173 = _RAND_2029[1:0];
  _RAND_2030 = {1{`RANDOM}};
  pht_7_174 = _RAND_2030[1:0];
  _RAND_2031 = {1{`RANDOM}};
  pht_7_175 = _RAND_2031[1:0];
  _RAND_2032 = {1{`RANDOM}};
  pht_7_176 = _RAND_2032[1:0];
  _RAND_2033 = {1{`RANDOM}};
  pht_7_177 = _RAND_2033[1:0];
  _RAND_2034 = {1{`RANDOM}};
  pht_7_178 = _RAND_2034[1:0];
  _RAND_2035 = {1{`RANDOM}};
  pht_7_179 = _RAND_2035[1:0];
  _RAND_2036 = {1{`RANDOM}};
  pht_7_180 = _RAND_2036[1:0];
  _RAND_2037 = {1{`RANDOM}};
  pht_7_181 = _RAND_2037[1:0];
  _RAND_2038 = {1{`RANDOM}};
  pht_7_182 = _RAND_2038[1:0];
  _RAND_2039 = {1{`RANDOM}};
  pht_7_183 = _RAND_2039[1:0];
  _RAND_2040 = {1{`RANDOM}};
  pht_7_184 = _RAND_2040[1:0];
  _RAND_2041 = {1{`RANDOM}};
  pht_7_185 = _RAND_2041[1:0];
  _RAND_2042 = {1{`RANDOM}};
  pht_7_186 = _RAND_2042[1:0];
  _RAND_2043 = {1{`RANDOM}};
  pht_7_187 = _RAND_2043[1:0];
  _RAND_2044 = {1{`RANDOM}};
  pht_7_188 = _RAND_2044[1:0];
  _RAND_2045 = {1{`RANDOM}};
  pht_7_189 = _RAND_2045[1:0];
  _RAND_2046 = {1{`RANDOM}};
  pht_7_190 = _RAND_2046[1:0];
  _RAND_2047 = {1{`RANDOM}};
  pht_7_191 = _RAND_2047[1:0];
  _RAND_2048 = {1{`RANDOM}};
  pht_7_192 = _RAND_2048[1:0];
  _RAND_2049 = {1{`RANDOM}};
  pht_7_193 = _RAND_2049[1:0];
  _RAND_2050 = {1{`RANDOM}};
  pht_7_194 = _RAND_2050[1:0];
  _RAND_2051 = {1{`RANDOM}};
  pht_7_195 = _RAND_2051[1:0];
  _RAND_2052 = {1{`RANDOM}};
  pht_7_196 = _RAND_2052[1:0];
  _RAND_2053 = {1{`RANDOM}};
  pht_7_197 = _RAND_2053[1:0];
  _RAND_2054 = {1{`RANDOM}};
  pht_7_198 = _RAND_2054[1:0];
  _RAND_2055 = {1{`RANDOM}};
  pht_7_199 = _RAND_2055[1:0];
  _RAND_2056 = {1{`RANDOM}};
  pht_7_200 = _RAND_2056[1:0];
  _RAND_2057 = {1{`RANDOM}};
  pht_7_201 = _RAND_2057[1:0];
  _RAND_2058 = {1{`RANDOM}};
  pht_7_202 = _RAND_2058[1:0];
  _RAND_2059 = {1{`RANDOM}};
  pht_7_203 = _RAND_2059[1:0];
  _RAND_2060 = {1{`RANDOM}};
  pht_7_204 = _RAND_2060[1:0];
  _RAND_2061 = {1{`RANDOM}};
  pht_7_205 = _RAND_2061[1:0];
  _RAND_2062 = {1{`RANDOM}};
  pht_7_206 = _RAND_2062[1:0];
  _RAND_2063 = {1{`RANDOM}};
  pht_7_207 = _RAND_2063[1:0];
  _RAND_2064 = {1{`RANDOM}};
  pht_7_208 = _RAND_2064[1:0];
  _RAND_2065 = {1{`RANDOM}};
  pht_7_209 = _RAND_2065[1:0];
  _RAND_2066 = {1{`RANDOM}};
  pht_7_210 = _RAND_2066[1:0];
  _RAND_2067 = {1{`RANDOM}};
  pht_7_211 = _RAND_2067[1:0];
  _RAND_2068 = {1{`RANDOM}};
  pht_7_212 = _RAND_2068[1:0];
  _RAND_2069 = {1{`RANDOM}};
  pht_7_213 = _RAND_2069[1:0];
  _RAND_2070 = {1{`RANDOM}};
  pht_7_214 = _RAND_2070[1:0];
  _RAND_2071 = {1{`RANDOM}};
  pht_7_215 = _RAND_2071[1:0];
  _RAND_2072 = {1{`RANDOM}};
  pht_7_216 = _RAND_2072[1:0];
  _RAND_2073 = {1{`RANDOM}};
  pht_7_217 = _RAND_2073[1:0];
  _RAND_2074 = {1{`RANDOM}};
  pht_7_218 = _RAND_2074[1:0];
  _RAND_2075 = {1{`RANDOM}};
  pht_7_219 = _RAND_2075[1:0];
  _RAND_2076 = {1{`RANDOM}};
  pht_7_220 = _RAND_2076[1:0];
  _RAND_2077 = {1{`RANDOM}};
  pht_7_221 = _RAND_2077[1:0];
  _RAND_2078 = {1{`RANDOM}};
  pht_7_222 = _RAND_2078[1:0];
  _RAND_2079 = {1{`RANDOM}};
  pht_7_223 = _RAND_2079[1:0];
  _RAND_2080 = {1{`RANDOM}};
  pht_7_224 = _RAND_2080[1:0];
  _RAND_2081 = {1{`RANDOM}};
  pht_7_225 = _RAND_2081[1:0];
  _RAND_2082 = {1{`RANDOM}};
  pht_7_226 = _RAND_2082[1:0];
  _RAND_2083 = {1{`RANDOM}};
  pht_7_227 = _RAND_2083[1:0];
  _RAND_2084 = {1{`RANDOM}};
  pht_7_228 = _RAND_2084[1:0];
  _RAND_2085 = {1{`RANDOM}};
  pht_7_229 = _RAND_2085[1:0];
  _RAND_2086 = {1{`RANDOM}};
  pht_7_230 = _RAND_2086[1:0];
  _RAND_2087 = {1{`RANDOM}};
  pht_7_231 = _RAND_2087[1:0];
  _RAND_2088 = {1{`RANDOM}};
  pht_7_232 = _RAND_2088[1:0];
  _RAND_2089 = {1{`RANDOM}};
  pht_7_233 = _RAND_2089[1:0];
  _RAND_2090 = {1{`RANDOM}};
  pht_7_234 = _RAND_2090[1:0];
  _RAND_2091 = {1{`RANDOM}};
  pht_7_235 = _RAND_2091[1:0];
  _RAND_2092 = {1{`RANDOM}};
  pht_7_236 = _RAND_2092[1:0];
  _RAND_2093 = {1{`RANDOM}};
  pht_7_237 = _RAND_2093[1:0];
  _RAND_2094 = {1{`RANDOM}};
  pht_7_238 = _RAND_2094[1:0];
  _RAND_2095 = {1{`RANDOM}};
  pht_7_239 = _RAND_2095[1:0];
  _RAND_2096 = {1{`RANDOM}};
  pht_7_240 = _RAND_2096[1:0];
  _RAND_2097 = {1{`RANDOM}};
  pht_7_241 = _RAND_2097[1:0];
  _RAND_2098 = {1{`RANDOM}};
  pht_7_242 = _RAND_2098[1:0];
  _RAND_2099 = {1{`RANDOM}};
  pht_7_243 = _RAND_2099[1:0];
  _RAND_2100 = {1{`RANDOM}};
  pht_7_244 = _RAND_2100[1:0];
  _RAND_2101 = {1{`RANDOM}};
  pht_7_245 = _RAND_2101[1:0];
  _RAND_2102 = {1{`RANDOM}};
  pht_7_246 = _RAND_2102[1:0];
  _RAND_2103 = {1{`RANDOM}};
  pht_7_247 = _RAND_2103[1:0];
  _RAND_2104 = {1{`RANDOM}};
  pht_7_248 = _RAND_2104[1:0];
  _RAND_2105 = {1{`RANDOM}};
  pht_7_249 = _RAND_2105[1:0];
  _RAND_2106 = {1{`RANDOM}};
  pht_7_250 = _RAND_2106[1:0];
  _RAND_2107 = {1{`RANDOM}};
  pht_7_251 = _RAND_2107[1:0];
  _RAND_2108 = {1{`RANDOM}};
  pht_7_252 = _RAND_2108[1:0];
  _RAND_2109 = {1{`RANDOM}};
  pht_7_253 = _RAND_2109[1:0];
  _RAND_2110 = {1{`RANDOM}};
  pht_7_254 = _RAND_2110[1:0];
  _RAND_2111 = {1{`RANDOM}};
  pht_7_255 = _RAND_2111[1:0];
  _RAND_2112 = {1{`RANDOM}};
  btb_0_valid = _RAND_2112[0:0];
  _RAND_2113 = {1{`RANDOM}};
  btb_0_tag = _RAND_2113[7:0];
  _RAND_2114 = {1{`RANDOM}};
  btb_0_target = _RAND_2114[31:0];
  _RAND_2115 = {1{`RANDOM}};
  btb_1_valid = _RAND_2115[0:0];
  _RAND_2116 = {1{`RANDOM}};
  btb_1_tag = _RAND_2116[7:0];
  _RAND_2117 = {1{`RANDOM}};
  btb_1_target = _RAND_2117[31:0];
  _RAND_2118 = {1{`RANDOM}};
  btb_2_valid = _RAND_2118[0:0];
  _RAND_2119 = {1{`RANDOM}};
  btb_2_tag = _RAND_2119[7:0];
  _RAND_2120 = {1{`RANDOM}};
  btb_2_target = _RAND_2120[31:0];
  _RAND_2121 = {1{`RANDOM}};
  btb_3_valid = _RAND_2121[0:0];
  _RAND_2122 = {1{`RANDOM}};
  btb_3_tag = _RAND_2122[7:0];
  _RAND_2123 = {1{`RANDOM}};
  btb_3_target = _RAND_2123[31:0];
  _RAND_2124 = {1{`RANDOM}};
  btb_4_valid = _RAND_2124[0:0];
  _RAND_2125 = {1{`RANDOM}};
  btb_4_tag = _RAND_2125[7:0];
  _RAND_2126 = {1{`RANDOM}};
  btb_4_target = _RAND_2126[31:0];
  _RAND_2127 = {1{`RANDOM}};
  btb_5_valid = _RAND_2127[0:0];
  _RAND_2128 = {1{`RANDOM}};
  btb_5_tag = _RAND_2128[7:0];
  _RAND_2129 = {1{`RANDOM}};
  btb_5_target = _RAND_2129[31:0];
  _RAND_2130 = {1{`RANDOM}};
  btb_6_valid = _RAND_2130[0:0];
  _RAND_2131 = {1{`RANDOM}};
  btb_6_tag = _RAND_2131[7:0];
  _RAND_2132 = {1{`RANDOM}};
  btb_6_target = _RAND_2132[31:0];
  _RAND_2133 = {1{`RANDOM}};
  btb_7_valid = _RAND_2133[0:0];
  _RAND_2134 = {1{`RANDOM}};
  btb_7_tag = _RAND_2134[7:0];
  _RAND_2135 = {1{`RANDOM}};
  btb_7_target = _RAND_2135[31:0];
  _RAND_2136 = {1{`RANDOM}};
  btb_8_valid = _RAND_2136[0:0];
  _RAND_2137 = {1{`RANDOM}};
  btb_8_tag = _RAND_2137[7:0];
  _RAND_2138 = {1{`RANDOM}};
  btb_8_target = _RAND_2138[31:0];
  _RAND_2139 = {1{`RANDOM}};
  btb_9_valid = _RAND_2139[0:0];
  _RAND_2140 = {1{`RANDOM}};
  btb_9_tag = _RAND_2140[7:0];
  _RAND_2141 = {1{`RANDOM}};
  btb_9_target = _RAND_2141[31:0];
  _RAND_2142 = {1{`RANDOM}};
  btb_10_valid = _RAND_2142[0:0];
  _RAND_2143 = {1{`RANDOM}};
  btb_10_tag = _RAND_2143[7:0];
  _RAND_2144 = {1{`RANDOM}};
  btb_10_target = _RAND_2144[31:0];
  _RAND_2145 = {1{`RANDOM}};
  btb_11_valid = _RAND_2145[0:0];
  _RAND_2146 = {1{`RANDOM}};
  btb_11_tag = _RAND_2146[7:0];
  _RAND_2147 = {1{`RANDOM}};
  btb_11_target = _RAND_2147[31:0];
  _RAND_2148 = {1{`RANDOM}};
  btb_12_valid = _RAND_2148[0:0];
  _RAND_2149 = {1{`RANDOM}};
  btb_12_tag = _RAND_2149[7:0];
  _RAND_2150 = {1{`RANDOM}};
  btb_12_target = _RAND_2150[31:0];
  _RAND_2151 = {1{`RANDOM}};
  btb_13_valid = _RAND_2151[0:0];
  _RAND_2152 = {1{`RANDOM}};
  btb_13_tag = _RAND_2152[7:0];
  _RAND_2153 = {1{`RANDOM}};
  btb_13_target = _RAND_2153[31:0];
  _RAND_2154 = {1{`RANDOM}};
  btb_14_valid = _RAND_2154[0:0];
  _RAND_2155 = {1{`RANDOM}};
  btb_14_tag = _RAND_2155[7:0];
  _RAND_2156 = {1{`RANDOM}};
  btb_14_target = _RAND_2156[31:0];
  _RAND_2157 = {1{`RANDOM}};
  btb_15_valid = _RAND_2157[0:0];
  _RAND_2158 = {1{`RANDOM}};
  btb_15_tag = _RAND_2158[7:0];
  _RAND_2159 = {1{`RANDOM}};
  btb_15_target = _RAND_2159[31:0];
  _RAND_2160 = {1{`RANDOM}};
  btb_16_valid = _RAND_2160[0:0];
  _RAND_2161 = {1{`RANDOM}};
  btb_16_tag = _RAND_2161[7:0];
  _RAND_2162 = {1{`RANDOM}};
  btb_16_target = _RAND_2162[31:0];
  _RAND_2163 = {1{`RANDOM}};
  btb_17_valid = _RAND_2163[0:0];
  _RAND_2164 = {1{`RANDOM}};
  btb_17_tag = _RAND_2164[7:0];
  _RAND_2165 = {1{`RANDOM}};
  btb_17_target = _RAND_2165[31:0];
  _RAND_2166 = {1{`RANDOM}};
  btb_18_valid = _RAND_2166[0:0];
  _RAND_2167 = {1{`RANDOM}};
  btb_18_tag = _RAND_2167[7:0];
  _RAND_2168 = {1{`RANDOM}};
  btb_18_target = _RAND_2168[31:0];
  _RAND_2169 = {1{`RANDOM}};
  btb_19_valid = _RAND_2169[0:0];
  _RAND_2170 = {1{`RANDOM}};
  btb_19_tag = _RAND_2170[7:0];
  _RAND_2171 = {1{`RANDOM}};
  btb_19_target = _RAND_2171[31:0];
  _RAND_2172 = {1{`RANDOM}};
  btb_20_valid = _RAND_2172[0:0];
  _RAND_2173 = {1{`RANDOM}};
  btb_20_tag = _RAND_2173[7:0];
  _RAND_2174 = {1{`RANDOM}};
  btb_20_target = _RAND_2174[31:0];
  _RAND_2175 = {1{`RANDOM}};
  btb_21_valid = _RAND_2175[0:0];
  _RAND_2176 = {1{`RANDOM}};
  btb_21_tag = _RAND_2176[7:0];
  _RAND_2177 = {1{`RANDOM}};
  btb_21_target = _RAND_2177[31:0];
  _RAND_2178 = {1{`RANDOM}};
  btb_22_valid = _RAND_2178[0:0];
  _RAND_2179 = {1{`RANDOM}};
  btb_22_tag = _RAND_2179[7:0];
  _RAND_2180 = {1{`RANDOM}};
  btb_22_target = _RAND_2180[31:0];
  _RAND_2181 = {1{`RANDOM}};
  btb_23_valid = _RAND_2181[0:0];
  _RAND_2182 = {1{`RANDOM}};
  btb_23_tag = _RAND_2182[7:0];
  _RAND_2183 = {1{`RANDOM}};
  btb_23_target = _RAND_2183[31:0];
  _RAND_2184 = {1{`RANDOM}};
  btb_24_valid = _RAND_2184[0:0];
  _RAND_2185 = {1{`RANDOM}};
  btb_24_tag = _RAND_2185[7:0];
  _RAND_2186 = {1{`RANDOM}};
  btb_24_target = _RAND_2186[31:0];
  _RAND_2187 = {1{`RANDOM}};
  btb_25_valid = _RAND_2187[0:0];
  _RAND_2188 = {1{`RANDOM}};
  btb_25_tag = _RAND_2188[7:0];
  _RAND_2189 = {1{`RANDOM}};
  btb_25_target = _RAND_2189[31:0];
  _RAND_2190 = {1{`RANDOM}};
  btb_26_valid = _RAND_2190[0:0];
  _RAND_2191 = {1{`RANDOM}};
  btb_26_tag = _RAND_2191[7:0];
  _RAND_2192 = {1{`RANDOM}};
  btb_26_target = _RAND_2192[31:0];
  _RAND_2193 = {1{`RANDOM}};
  btb_27_valid = _RAND_2193[0:0];
  _RAND_2194 = {1{`RANDOM}};
  btb_27_tag = _RAND_2194[7:0];
  _RAND_2195 = {1{`RANDOM}};
  btb_27_target = _RAND_2195[31:0];
  _RAND_2196 = {1{`RANDOM}};
  btb_28_valid = _RAND_2196[0:0];
  _RAND_2197 = {1{`RANDOM}};
  btb_28_tag = _RAND_2197[7:0];
  _RAND_2198 = {1{`RANDOM}};
  btb_28_target = _RAND_2198[31:0];
  _RAND_2199 = {1{`RANDOM}};
  btb_29_valid = _RAND_2199[0:0];
  _RAND_2200 = {1{`RANDOM}};
  btb_29_tag = _RAND_2200[7:0];
  _RAND_2201 = {1{`RANDOM}};
  btb_29_target = _RAND_2201[31:0];
  _RAND_2202 = {1{`RANDOM}};
  btb_30_valid = _RAND_2202[0:0];
  _RAND_2203 = {1{`RANDOM}};
  btb_30_tag = _RAND_2203[7:0];
  _RAND_2204 = {1{`RANDOM}};
  btb_30_target = _RAND_2204[31:0];
  _RAND_2205 = {1{`RANDOM}};
  btb_31_valid = _RAND_2205[0:0];
  _RAND_2206 = {1{`RANDOM}};
  btb_31_tag = _RAND_2206[7:0];
  _RAND_2207 = {1{`RANDOM}};
  btb_31_target = _RAND_2207[31:0];
  _RAND_2208 = {1{`RANDOM}};
  btb_32_valid = _RAND_2208[0:0];
  _RAND_2209 = {1{`RANDOM}};
  btb_32_tag = _RAND_2209[7:0];
  _RAND_2210 = {1{`RANDOM}};
  btb_32_target = _RAND_2210[31:0];
  _RAND_2211 = {1{`RANDOM}};
  btb_33_valid = _RAND_2211[0:0];
  _RAND_2212 = {1{`RANDOM}};
  btb_33_tag = _RAND_2212[7:0];
  _RAND_2213 = {1{`RANDOM}};
  btb_33_target = _RAND_2213[31:0];
  _RAND_2214 = {1{`RANDOM}};
  btb_34_valid = _RAND_2214[0:0];
  _RAND_2215 = {1{`RANDOM}};
  btb_34_tag = _RAND_2215[7:0];
  _RAND_2216 = {1{`RANDOM}};
  btb_34_target = _RAND_2216[31:0];
  _RAND_2217 = {1{`RANDOM}};
  btb_35_valid = _RAND_2217[0:0];
  _RAND_2218 = {1{`RANDOM}};
  btb_35_tag = _RAND_2218[7:0];
  _RAND_2219 = {1{`RANDOM}};
  btb_35_target = _RAND_2219[31:0];
  _RAND_2220 = {1{`RANDOM}};
  btb_36_valid = _RAND_2220[0:0];
  _RAND_2221 = {1{`RANDOM}};
  btb_36_tag = _RAND_2221[7:0];
  _RAND_2222 = {1{`RANDOM}};
  btb_36_target = _RAND_2222[31:0];
  _RAND_2223 = {1{`RANDOM}};
  btb_37_valid = _RAND_2223[0:0];
  _RAND_2224 = {1{`RANDOM}};
  btb_37_tag = _RAND_2224[7:0];
  _RAND_2225 = {1{`RANDOM}};
  btb_37_target = _RAND_2225[31:0];
  _RAND_2226 = {1{`RANDOM}};
  btb_38_valid = _RAND_2226[0:0];
  _RAND_2227 = {1{`RANDOM}};
  btb_38_tag = _RAND_2227[7:0];
  _RAND_2228 = {1{`RANDOM}};
  btb_38_target = _RAND_2228[31:0];
  _RAND_2229 = {1{`RANDOM}};
  btb_39_valid = _RAND_2229[0:0];
  _RAND_2230 = {1{`RANDOM}};
  btb_39_tag = _RAND_2230[7:0];
  _RAND_2231 = {1{`RANDOM}};
  btb_39_target = _RAND_2231[31:0];
  _RAND_2232 = {1{`RANDOM}};
  btb_40_valid = _RAND_2232[0:0];
  _RAND_2233 = {1{`RANDOM}};
  btb_40_tag = _RAND_2233[7:0];
  _RAND_2234 = {1{`RANDOM}};
  btb_40_target = _RAND_2234[31:0];
  _RAND_2235 = {1{`RANDOM}};
  btb_41_valid = _RAND_2235[0:0];
  _RAND_2236 = {1{`RANDOM}};
  btb_41_tag = _RAND_2236[7:0];
  _RAND_2237 = {1{`RANDOM}};
  btb_41_target = _RAND_2237[31:0];
  _RAND_2238 = {1{`RANDOM}};
  btb_42_valid = _RAND_2238[0:0];
  _RAND_2239 = {1{`RANDOM}};
  btb_42_tag = _RAND_2239[7:0];
  _RAND_2240 = {1{`RANDOM}};
  btb_42_target = _RAND_2240[31:0];
  _RAND_2241 = {1{`RANDOM}};
  btb_43_valid = _RAND_2241[0:0];
  _RAND_2242 = {1{`RANDOM}};
  btb_43_tag = _RAND_2242[7:0];
  _RAND_2243 = {1{`RANDOM}};
  btb_43_target = _RAND_2243[31:0];
  _RAND_2244 = {1{`RANDOM}};
  btb_44_valid = _RAND_2244[0:0];
  _RAND_2245 = {1{`RANDOM}};
  btb_44_tag = _RAND_2245[7:0];
  _RAND_2246 = {1{`RANDOM}};
  btb_44_target = _RAND_2246[31:0];
  _RAND_2247 = {1{`RANDOM}};
  btb_45_valid = _RAND_2247[0:0];
  _RAND_2248 = {1{`RANDOM}};
  btb_45_tag = _RAND_2248[7:0];
  _RAND_2249 = {1{`RANDOM}};
  btb_45_target = _RAND_2249[31:0];
  _RAND_2250 = {1{`RANDOM}};
  btb_46_valid = _RAND_2250[0:0];
  _RAND_2251 = {1{`RANDOM}};
  btb_46_tag = _RAND_2251[7:0];
  _RAND_2252 = {1{`RANDOM}};
  btb_46_target = _RAND_2252[31:0];
  _RAND_2253 = {1{`RANDOM}};
  btb_47_valid = _RAND_2253[0:0];
  _RAND_2254 = {1{`RANDOM}};
  btb_47_tag = _RAND_2254[7:0];
  _RAND_2255 = {1{`RANDOM}};
  btb_47_target = _RAND_2255[31:0];
  _RAND_2256 = {1{`RANDOM}};
  btb_48_valid = _RAND_2256[0:0];
  _RAND_2257 = {1{`RANDOM}};
  btb_48_tag = _RAND_2257[7:0];
  _RAND_2258 = {1{`RANDOM}};
  btb_48_target = _RAND_2258[31:0];
  _RAND_2259 = {1{`RANDOM}};
  btb_49_valid = _RAND_2259[0:0];
  _RAND_2260 = {1{`RANDOM}};
  btb_49_tag = _RAND_2260[7:0];
  _RAND_2261 = {1{`RANDOM}};
  btb_49_target = _RAND_2261[31:0];
  _RAND_2262 = {1{`RANDOM}};
  btb_50_valid = _RAND_2262[0:0];
  _RAND_2263 = {1{`RANDOM}};
  btb_50_tag = _RAND_2263[7:0];
  _RAND_2264 = {1{`RANDOM}};
  btb_50_target = _RAND_2264[31:0];
  _RAND_2265 = {1{`RANDOM}};
  btb_51_valid = _RAND_2265[0:0];
  _RAND_2266 = {1{`RANDOM}};
  btb_51_tag = _RAND_2266[7:0];
  _RAND_2267 = {1{`RANDOM}};
  btb_51_target = _RAND_2267[31:0];
  _RAND_2268 = {1{`RANDOM}};
  btb_52_valid = _RAND_2268[0:0];
  _RAND_2269 = {1{`RANDOM}};
  btb_52_tag = _RAND_2269[7:0];
  _RAND_2270 = {1{`RANDOM}};
  btb_52_target = _RAND_2270[31:0];
  _RAND_2271 = {1{`RANDOM}};
  btb_53_valid = _RAND_2271[0:0];
  _RAND_2272 = {1{`RANDOM}};
  btb_53_tag = _RAND_2272[7:0];
  _RAND_2273 = {1{`RANDOM}};
  btb_53_target = _RAND_2273[31:0];
  _RAND_2274 = {1{`RANDOM}};
  btb_54_valid = _RAND_2274[0:0];
  _RAND_2275 = {1{`RANDOM}};
  btb_54_tag = _RAND_2275[7:0];
  _RAND_2276 = {1{`RANDOM}};
  btb_54_target = _RAND_2276[31:0];
  _RAND_2277 = {1{`RANDOM}};
  btb_55_valid = _RAND_2277[0:0];
  _RAND_2278 = {1{`RANDOM}};
  btb_55_tag = _RAND_2278[7:0];
  _RAND_2279 = {1{`RANDOM}};
  btb_55_target = _RAND_2279[31:0];
  _RAND_2280 = {1{`RANDOM}};
  btb_56_valid = _RAND_2280[0:0];
  _RAND_2281 = {1{`RANDOM}};
  btb_56_tag = _RAND_2281[7:0];
  _RAND_2282 = {1{`RANDOM}};
  btb_56_target = _RAND_2282[31:0];
  _RAND_2283 = {1{`RANDOM}};
  btb_57_valid = _RAND_2283[0:0];
  _RAND_2284 = {1{`RANDOM}};
  btb_57_tag = _RAND_2284[7:0];
  _RAND_2285 = {1{`RANDOM}};
  btb_57_target = _RAND_2285[31:0];
  _RAND_2286 = {1{`RANDOM}};
  btb_58_valid = _RAND_2286[0:0];
  _RAND_2287 = {1{`RANDOM}};
  btb_58_tag = _RAND_2287[7:0];
  _RAND_2288 = {1{`RANDOM}};
  btb_58_target = _RAND_2288[31:0];
  _RAND_2289 = {1{`RANDOM}};
  btb_59_valid = _RAND_2289[0:0];
  _RAND_2290 = {1{`RANDOM}};
  btb_59_tag = _RAND_2290[7:0];
  _RAND_2291 = {1{`RANDOM}};
  btb_59_target = _RAND_2291[31:0];
  _RAND_2292 = {1{`RANDOM}};
  btb_60_valid = _RAND_2292[0:0];
  _RAND_2293 = {1{`RANDOM}};
  btb_60_tag = _RAND_2293[7:0];
  _RAND_2294 = {1{`RANDOM}};
  btb_60_target = _RAND_2294[31:0];
  _RAND_2295 = {1{`RANDOM}};
  btb_61_valid = _RAND_2295[0:0];
  _RAND_2296 = {1{`RANDOM}};
  btb_61_tag = _RAND_2296[7:0];
  _RAND_2297 = {1{`RANDOM}};
  btb_61_target = _RAND_2297[31:0];
  _RAND_2298 = {1{`RANDOM}};
  btb_62_valid = _RAND_2298[0:0];
  _RAND_2299 = {1{`RANDOM}};
  btb_62_tag = _RAND_2299[7:0];
  _RAND_2300 = {1{`RANDOM}};
  btb_62_target = _RAND_2300[31:0];
  _RAND_2301 = {1{`RANDOM}};
  btb_63_valid = _RAND_2301[0:0];
  _RAND_2302 = {1{`RANDOM}};
  btb_63_tag = _RAND_2302[7:0];
  _RAND_2303 = {1{`RANDOM}};
  btb_63_target = _RAND_2303[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InstFetch(
  input         clock,
  input         reset,
  output        io_imem_inst_valid,
  input         io_imem_inst_ready,
  output [31:0] io_imem_inst_addr,
  input  [31:0] io_imem_inst_read,
  input         io_jmp_packet_valid,
  input  [31:0] io_jmp_packet_inst_pc,
  input         io_jmp_packet_jmp,
  input  [31:0] io_jmp_packet_jmp_pc,
  input         io_jmp_packet_mis,
  input         io_stall,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_bp_taken,
  output [31:0] io_out_bp_targer
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  bp_clock; // @[InstFetch.scala 20:18]
  wire  bp_reset; // @[InstFetch.scala 20:18]
  wire [31:0] bp_io_pc; // @[InstFetch.scala 20:18]
  wire  bp_io_is_br; // @[InstFetch.scala 20:18]
  wire  bp_io_jmp_packet_valid; // @[InstFetch.scala 20:18]
  wire [31:0] bp_io_jmp_packet_inst_pc; // @[InstFetch.scala 20:18]
  wire  bp_io_jmp_packet_jmp; // @[InstFetch.scala 20:18]
  wire [31:0] bp_io_jmp_packet_jmp_pc; // @[InstFetch.scala 20:18]
  wire  bp_io_jmp_packet_mis; // @[InstFetch.scala 20:18]
  wire  bp_io_pred_br; // @[InstFetch.scala 20:18]
  wire [31:0] bp_io_pred_pc; // @[InstFetch.scala 20:18]
  reg [31:0] pc; // @[InstFetch.scala 18:19]
  reg [31:0] inst; // @[InstFetch.scala 19:21]
  reg  reg_mis; // @[InstFetch.scala 24:24]
  reg [31:0] mis_pc; // @[InstFetch.scala 25:24]
  wire [31:0] _mis_pc_T_1 = io_jmp_packet_inst_pc + 32'h4; // @[InstFetch.scala 28:83]
  wire  _T = ~io_jmp_packet_mis; // @[InstFetch.scala 29:38]
  wire  _GEN_0 = io_imem_inst_ready & ~io_jmp_packet_mis ? 1'h0 : reg_mis; // @[InstFetch.scala 29:44 InstFetch.scala 30:13 InstFetch.scala 24:24]
  wire  _GEN_2 = io_jmp_packet_mis | _GEN_0; // @[InstFetch.scala 26:14 InstFetch.scala 27:13]
  wire  _io_imem_inst_valid_T = ~io_stall; // @[InstFetch.scala 36:25]
  wire [31:0] _bp_io_is_br_T = inst & 32'h7f; // @[InstFetch.scala 44:24]
  wire [31:0] _bp_io_is_br_T_2 = inst & 32'h707f; // @[InstFetch.scala 44:55]
  wire  _bp_io_is_br_T_6 = 32'h63 == _bp_io_is_br_T_2; // @[InstFetch.scala 45:24]
  wire  _bp_io_is_br_T_7 = 32'h6f == _bp_io_is_br_T | 32'h67 == _bp_io_is_br_T_2 | _bp_io_is_br_T_6; // @[InstFetch.scala 44:78]
  wire  _bp_io_is_br_T_12 = 32'h4063 == _bp_io_is_br_T_2; // @[InstFetch.scala 46:24]
  wire  _bp_io_is_br_T_13 = _bp_io_is_br_T_7 | 32'h1063 == _bp_io_is_br_T_2 | _bp_io_is_br_T_12; // @[InstFetch.scala 45:78]
  wire  _bp_io_is_br_T_18 = 32'h5063 == _bp_io_is_br_T_2; // @[InstFetch.scala 47:24]
  wire  _bp_io_is_br_T_19 = _bp_io_is_br_T_13 | 32'h6063 == _bp_io_is_br_T_2 | _bp_io_is_br_T_18; // @[InstFetch.scala 46:78]
  wire  _T_3 = io_imem_inst_ready & _io_imem_inst_valid_T; // @[InstFetch.scala 51:19]
  reg  if_stall; // @[InstFetch.scala 57:25]
  reg  if_valid; // @[InstFetch.scala 58:25]
  wire  _GEN_6 = _io_imem_inst_valid_T ? 1'h0 : if_stall; // @[InstFetch.scala 61:23 InstFetch.scala 62:14 InstFetch.scala 57:25]
  wire  _GEN_7 = if_valid & io_stall | _GEN_6; // @[InstFetch.scala 59:28 InstFetch.scala 60:14]
  wire  _if_pc_T = io_jmp_packet_mis | reg_mis; // @[InstFetch.scala 70:25]
  BrPredictor bp ( // @[InstFetch.scala 20:18]
    .clock(bp_clock),
    .reset(bp_reset),
    .io_pc(bp_io_pc),
    .io_is_br(bp_io_is_br),
    .io_jmp_packet_valid(bp_io_jmp_packet_valid),
    .io_jmp_packet_inst_pc(bp_io_jmp_packet_inst_pc),
    .io_jmp_packet_jmp(bp_io_jmp_packet_jmp),
    .io_jmp_packet_jmp_pc(bp_io_jmp_packet_jmp_pc),
    .io_jmp_packet_mis(bp_io_jmp_packet_mis),
    .io_pred_br(bp_io_pred_br),
    .io_pred_pc(bp_io_pred_pc)
  );
  assign io_imem_inst_valid = ~io_stall; // @[InstFetch.scala 36:25]
  assign io_imem_inst_addr = reg_mis ? mis_pc : bp_io_pred_pc; // @[InstFetch.scala 34:16]
  assign io_out_valid = (if_valid | if_stall) & _T & ~reg_mis; // @[InstFetch.scala 73:55]
  assign io_out_pc = io_jmp_packet_mis | reg_mis ? 32'h0 : pc; // @[InstFetch.scala 70:20]
  assign io_out_inst = _if_pc_T ? 32'h0 : inst; // @[InstFetch.scala 71:20]
  assign io_out_bp_taken = bp_io_pred_br; // @[InstFetch.scala 89:21]
  assign io_out_bp_targer = bp_io_pred_pc; // @[InstFetch.scala 90:21]
  assign bp_clock = clock;
  assign bp_reset = reset;
  assign bp_io_pc = pc; // @[InstFetch.scala 42:12]
  assign bp_io_is_br = _bp_io_is_br_T_19 | 32'h7063 == _bp_io_is_br_T_2; // @[InstFetch.scala 47:46]
  assign bp_io_jmp_packet_valid = io_jmp_packet_valid; // @[InstFetch.scala 48:20]
  assign bp_io_jmp_packet_inst_pc = io_jmp_packet_inst_pc; // @[InstFetch.scala 48:20]
  assign bp_io_jmp_packet_jmp = io_jmp_packet_jmp; // @[InstFetch.scala 48:20]
  assign bp_io_jmp_packet_jmp_pc = io_jmp_packet_jmp_pc; // @[InstFetch.scala 48:20]
  assign bp_io_jmp_packet_mis = io_jmp_packet_mis; // @[InstFetch.scala 48:20]
  always @(posedge clock) begin
    if (reset) begin // @[InstFetch.scala 18:19]
      pc <= 32'h7ffffffc; // @[InstFetch.scala 18:19]
    end else if (io_imem_inst_ready & _io_imem_inst_valid_T) begin // @[InstFetch.scala 51:30]
      if (reg_mis) begin // @[InstFetch.scala 34:16]
        pc <= mis_pc;
      end else begin
        pc <= bp_io_pred_pc;
      end
    end
    if (reset) begin // @[InstFetch.scala 19:21]
      inst <= 32'h0; // @[InstFetch.scala 19:21]
    end else if (io_imem_inst_ready & _io_imem_inst_valid_T) begin // @[InstFetch.scala 51:30]
      inst <= io_imem_inst_read; // @[InstFetch.scala 53:11]
    end
    if (reset) begin // @[InstFetch.scala 24:24]
      reg_mis <= 1'h0; // @[InstFetch.scala 24:24]
    end else begin
      reg_mis <= _GEN_2;
    end
    if (reset) begin // @[InstFetch.scala 25:24]
      mis_pc <= 32'h0; // @[InstFetch.scala 25:24]
    end else if (io_jmp_packet_mis) begin // @[InstFetch.scala 26:14]
      if (io_jmp_packet_jmp) begin // @[InstFetch.scala 28:19]
        mis_pc <= io_jmp_packet_jmp_pc;
      end else begin
        mis_pc <= _mis_pc_T_1;
      end
    end else if (io_imem_inst_ready & ~io_jmp_packet_mis) begin // @[InstFetch.scala 29:44]
      mis_pc <= 32'h0; // @[InstFetch.scala 31:13]
    end
    if (reset) begin // @[InstFetch.scala 57:25]
      if_stall <= 1'h0; // @[InstFetch.scala 57:25]
    end else begin
      if_stall <= _GEN_7;
    end
    if (reset) begin // @[InstFetch.scala 58:25]
      if_valid <= 1'h0; // @[InstFetch.scala 58:25]
    end else begin
      if_valid <= _T_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  inst = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_mis = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  mis_pc = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  if_stall = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  if_valid = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelineReg(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_wen,
  input  [4:0]  io_in_wdest,
  input  [63:0] io_in_wdata,
  input  [63:0] io_in_op1,
  input  [63:0] io_in_op2,
  input         io_in_typew,
  input  [63:0] io_in_wmem,
  input  [31:0] io_in_mem_addr,
  input  [11:0] io_in_aluop,
  input  [6:0]  io_in_loadop,
  input  [3:0]  io_in_storeop,
  input  [3:0]  io_in_sysop,
  input         io_in_bp_taken,
  input  [31:0] io_in_bp_targer,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_wen,
  output [4:0]  io_out_wdest,
  output [63:0] io_out_wdata,
  output [63:0] io_out_op1,
  output [63:0] io_out_op2,
  output        io_out_typew,
  output [63:0] io_out_wmem,
  output [31:0] io_out_mem_addr,
  output [11:0] io_out_aluop,
  output [6:0]  io_out_loadop,
  output [3:0]  io_out_storeop,
  output [3:0]  io_out_sysop,
  output        io_out_bp_taken,
  output [31:0] io_out_bp_targer,
  input         io_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg  reg_valid; // @[PipelineReg.scala 57:20]
  reg [31:0] reg_pc; // @[PipelineReg.scala 57:20]
  reg [31:0] reg_inst; // @[PipelineReg.scala 57:20]
  reg  reg_wen; // @[PipelineReg.scala 57:20]
  reg [4:0] reg_wdest; // @[PipelineReg.scala 57:20]
  reg [63:0] reg_wdata; // @[PipelineReg.scala 57:20]
  reg [63:0] reg_op1; // @[PipelineReg.scala 57:20]
  reg [63:0] reg_op2; // @[PipelineReg.scala 57:20]
  reg  reg_typew; // @[PipelineReg.scala 57:20]
  reg [63:0] reg_wmem; // @[PipelineReg.scala 57:20]
  reg [31:0] reg_mem_addr; // @[PipelineReg.scala 57:20]
  reg [11:0] reg_aluop; // @[PipelineReg.scala 57:20]
  reg [6:0] reg_loadop; // @[PipelineReg.scala 57:20]
  reg [3:0] reg_storeop; // @[PipelineReg.scala 57:20]
  reg [3:0] reg_sysop; // @[PipelineReg.scala 57:20]
  reg  reg_bp_taken; // @[PipelineReg.scala 57:20]
  reg [31:0] reg_bp_targer; // @[PipelineReg.scala 57:20]
  wire  _T = ~io_stall; // @[PipelineReg.scala 59:21]
  assign io_out_valid = reg_valid; // @[PipelineReg.scala 65:10]
  assign io_out_pc = reg_pc; // @[PipelineReg.scala 65:10]
  assign io_out_inst = reg_inst; // @[PipelineReg.scala 65:10]
  assign io_out_wen = reg_wen; // @[PipelineReg.scala 65:10]
  assign io_out_wdest = reg_wdest; // @[PipelineReg.scala 65:10]
  assign io_out_wdata = reg_wdata; // @[PipelineReg.scala 65:10]
  assign io_out_op1 = reg_op1; // @[PipelineReg.scala 65:10]
  assign io_out_op2 = reg_op2; // @[PipelineReg.scala 65:10]
  assign io_out_typew = reg_typew; // @[PipelineReg.scala 65:10]
  assign io_out_wmem = reg_wmem; // @[PipelineReg.scala 65:10]
  assign io_out_mem_addr = reg_mem_addr; // @[PipelineReg.scala 65:10]
  assign io_out_aluop = reg_aluop; // @[PipelineReg.scala 65:10]
  assign io_out_loadop = reg_loadop; // @[PipelineReg.scala 65:10]
  assign io_out_storeop = reg_storeop; // @[PipelineReg.scala 65:10]
  assign io_out_sysop = reg_sysop; // @[PipelineReg.scala 65:10]
  assign io_out_bp_taken = reg_bp_taken; // @[PipelineReg.scala 65:10]
  assign io_out_bp_targer = reg_bp_targer; // @[PipelineReg.scala 65:10]
  always @(posedge clock) begin
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_valid <= 1'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_valid <= io_in_valid; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_pc <= 32'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_pc <= io_in_pc; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_inst <= 32'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_inst <= io_in_inst; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_wen <= 1'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_wen <= io_in_wen; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_wdest <= 5'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_wdest <= io_in_wdest; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_wdata <= 64'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_wdata <= io_in_wdata; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_op1 <= 64'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_op1 <= io_in_op1; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_op2 <= 64'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_op2 <= io_in_op2; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_typew <= 1'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_typew <= io_in_typew; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_wmem <= 64'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_wmem <= io_in_wmem; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_mem_addr <= 32'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_mem_addr <= io_in_mem_addr; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_aluop <= 12'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_aluop <= io_in_aluop; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_loadop <= 7'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_loadop <= io_in_loadop; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_storeop <= 4'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_storeop <= io_in_storeop; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_sysop <= 4'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_sysop <= io_in_sysop; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_bp_taken <= 1'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_bp_taken <= io_in_bp_taken; // @[PipelineReg.scala 62:9]
    end
    if (reset) begin // @[PipelineReg.scala 57:20]
      reg_bp_targer <= 32'h0; // @[PipelineReg.scala 57:20]
    end else if (_T) begin // @[PipelineReg.scala 61:27]
      reg_bp_targer <= io_in_bp_targer; // @[PipelineReg.scala 62:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_wen = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reg_wdest = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  reg_wdata = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  reg_op1 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  reg_op2 = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  reg_typew = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  reg_wmem = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  reg_mem_addr = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_aluop = _RAND_11[11:0];
  _RAND_12 = {1{`RANDOM}};
  reg_loadop = _RAND_12[6:0];
  _RAND_13 = {1{`RANDOM}};
  reg_storeop = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  reg_sysop = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  reg_bp_taken = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  reg_bp_targer = _RAND_16[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Ctrl(
  input  [10:0] io_redirectop,
  input  [31:0] io_pc,
  input  [31:0] io_imm_i,
  input  [31:0] io_imm_j,
  input  [31:0] io_imm_b,
  input  [63:0] io_rs1_value,
  input  [63:0] io_rs2_value,
  input  [63:0] io_mtvec,
  input  [63:0] io_mepc,
  output        io_jmp,
  output [63:0] io_target
);
  wire  _io_jmp_T_2 = io_redirectop == 11'h2; // @[Ctrl.scala 32:29]
  wire  _io_jmp_T_4 = io_redirectop == 11'h4 | _io_jmp_T_2; // @[Ctrl.scala 31:66]
  wire  _io_jmp_T_5 = io_redirectop == 11'h1; // @[Ctrl.scala 33:29]
  wire  _io_jmp_T_7 = _io_jmp_T_4 | _io_jmp_T_5; // @[Ctrl.scala 32:66]
  wire  _io_jmp_T_8 = io_redirectop == 11'h10; // @[Ctrl.scala 34:29]
  wire  _io_jmp_T_10 = _io_jmp_T_7 | _io_jmp_T_8; // @[Ctrl.scala 33:66]
  wire  _io_jmp_T_11 = io_redirectop == 11'h8; // @[Ctrl.scala 35:29]
  wire  _io_jmp_T_13 = _io_jmp_T_10 | _io_jmp_T_11; // @[Ctrl.scala 34:66]
  wire  _io_jmp_T_16 = io_redirectop == 11'h400 & io_rs1_value == io_rs2_value; // @[Ctrl.scala 36:55]
  wire  _io_jmp_T_17 = _io_jmp_T_13 | _io_jmp_T_16; // @[Ctrl.scala 35:66]
  wire  _io_jmp_T_20 = io_redirectop == 11'h200 & io_rs1_value != io_rs2_value; // @[Ctrl.scala 37:55]
  wire  _io_jmp_T_21 = _io_jmp_T_17 | _io_jmp_T_20; // @[Ctrl.scala 36:83]
  wire  _io_jmp_T_26 = io_redirectop == 11'h100 & $signed(io_rs1_value) < $signed(io_rs2_value); // @[Ctrl.scala 38:55]
  wire  _io_jmp_T_27 = _io_jmp_T_21 | _io_jmp_T_26; // @[Ctrl.scala 37:83]
  wire  _io_jmp_T_32 = io_redirectop == 11'h80 & $signed(io_rs1_value) >= $signed(io_rs2_value); // @[Ctrl.scala 39:55]
  wire  _io_jmp_T_33 = _io_jmp_T_27 | _io_jmp_T_32; // @[Ctrl.scala 38:100]
  wire  _io_jmp_T_36 = io_redirectop == 11'h40 & io_rs1_value < io_rs2_value; // @[Ctrl.scala 40:55]
  wire  _io_jmp_T_37 = _io_jmp_T_33 | _io_jmp_T_36; // @[Ctrl.scala 39:100]
  wire  _io_jmp_T_40 = io_redirectop == 11'h20 & io_rs1_value >= io_rs2_value; // @[Ctrl.scala 41:55]
  wire [29:0] io_target_hi = io_mtvec[31:2]; // @[Ctrl.scala 44:53]
  wire [31:0] _io_target_T = {io_target_hi,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] _io_target_T_4 = io_pc + io_imm_j; // @[Ctrl.scala 47:48]
  wire [63:0] _GEN_0 = {{32'd0}, io_imm_i}; // @[Ctrl.scala 48:55]
  wire [63:0] _io_target_T_6 = io_rs1_value + _GEN_0; // @[Ctrl.scala 48:55]
  wire [31:0] _io_target_T_8 = io_pc + io_imm_b; // @[Ctrl.scala 49:48]
  wire [31:0] _io_target_T_20 = 11'h4 == io_redirectop ? _io_target_T : 32'h0; // @[Mux.scala 80:57]
  wire [31:0] _io_target_T_22 = 11'h2 == io_redirectop ? io_mepc[31:0] : _io_target_T_20; // @[Mux.scala 80:57]
  wire [31:0] _io_target_T_24 = 11'h1 == io_redirectop ? _io_target_T : _io_target_T_22; // @[Mux.scala 80:57]
  wire [31:0] _io_target_T_26 = 11'h10 == io_redirectop ? _io_target_T_4 : _io_target_T_24; // @[Mux.scala 80:57]
  wire [63:0] _io_target_T_28 = 11'h8 == io_redirectop ? _io_target_T_6 : {{32'd0}, _io_target_T_26}; // @[Mux.scala 80:57]
  wire [63:0] _io_target_T_30 = 11'h400 == io_redirectop ? {{32'd0}, _io_target_T_8} : _io_target_T_28; // @[Mux.scala 80:57]
  wire [63:0] _io_target_T_32 = 11'h200 == io_redirectop ? {{32'd0}, _io_target_T_8} : _io_target_T_30; // @[Mux.scala 80:57]
  wire [63:0] _io_target_T_34 = 11'h100 == io_redirectop ? {{32'd0}, _io_target_T_8} : _io_target_T_32; // @[Mux.scala 80:57]
  wire [63:0] _io_target_T_36 = 11'h80 == io_redirectop ? {{32'd0}, _io_target_T_8} : _io_target_T_34; // @[Mux.scala 80:57]
  wire [63:0] _io_target_T_38 = 11'h40 == io_redirectop ? {{32'd0}, _io_target_T_8} : _io_target_T_36; // @[Mux.scala 80:57]
  assign io_jmp = _io_jmp_T_37 | _io_jmp_T_40; // @[Ctrl.scala 40:100]
  assign io_target = 11'h20 == io_redirectop ? {{32'd0}, _io_target_T_8} : _io_target_T_38; // @[Mux.scala 80:57]
endmodule
module Decode(
  output [4:0]  io_rs1_addr,
  output [4:0]  io_rs2_addr,
  input  [63:0] io_rs1_data,
  input  [63:0] io_rs2_data,
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_bp_taken,
  input  [31:0] io_in_bp_targer,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_wen,
  output [4:0]  io_out_wdest,
  output [63:0] io_out_op1,
  output [63:0] io_out_op2,
  output        io_out_typew,
  output [63:0] io_out_wmem,
  output [11:0] io_out_aluop,
  output [6:0]  io_out_loadop,
  output [3:0]  io_out_storeop,
  output [3:0]  io_out_sysop,
  output        io_jmp_packet_valid,
  output [31:0] io_jmp_packet_inst_pc,
  output        io_jmp_packet_jmp,
  output [31:0] io_jmp_packet_jmp_pc,
  output        io_jmp_packet_mis,
  input         io_stall,
  input  [63:0] io_mtvec,
  input  [63:0] io_mepc,
  input         io_time_int,
  input  [4:0]  io_ex_wdest,
  input  [4:0]  io_wb_wdest,
  input  [63:0] io_ex_result,
  input  [63:0] io_wb_result
);
  wire [10:0] ctrl_io_redirectop; // @[Decode.scala 217:20]
  wire [31:0] ctrl_io_pc; // @[Decode.scala 217:20]
  wire [31:0] ctrl_io_imm_i; // @[Decode.scala 217:20]
  wire [31:0] ctrl_io_imm_j; // @[Decode.scala 217:20]
  wire [31:0] ctrl_io_imm_b; // @[Decode.scala 217:20]
  wire [63:0] ctrl_io_rs1_value; // @[Decode.scala 217:20]
  wire [63:0] ctrl_io_rs2_value; // @[Decode.scala 217:20]
  wire [63:0] ctrl_io_mtvec; // @[Decode.scala 217:20]
  wire [63:0] ctrl_io_mepc; // @[Decode.scala 217:20]
  wire  ctrl_io_jmp; // @[Decode.scala 217:20]
  wire [63:0] ctrl_io_target; // @[Decode.scala 217:20]
  wire [31:0] _addi_T = io_in_inst & 32'h707f; // @[Decode.scala 39:22]
  wire  addi = 32'h13 == _addi_T; // @[Decode.scala 39:22]
  wire  andi = 32'h7013 == _addi_T; // @[Decode.scala 40:22]
  wire  xori = 32'h4013 == _addi_T; // @[Decode.scala 41:22]
  wire  ori = 32'h6013 == _addi_T; // @[Decode.scala 42:22]
  wire [31:0] _slli_T = io_in_inst & 32'hfc00707f; // @[Decode.scala 43:22]
  wire  slli = 32'h1013 == _slli_T; // @[Decode.scala 43:22]
  wire  srli = 32'h5013 == _slli_T; // @[Decode.scala 44:22]
  wire  srai = 32'h40005013 == _slli_T; // @[Decode.scala 45:22]
  wire  slti = 32'h2013 == _addi_T; // @[Decode.scala 46:22]
  wire  sltiu = 32'h3013 == _addi_T; // @[Decode.scala 47:22]
  wire  addiw = 32'h1b == _addi_T; // @[Decode.scala 48:22]
  wire [31:0] _slliw_T = io_in_inst & 32'hfe00707f; // @[Decode.scala 49:22]
  wire  slliw = 32'h101b == _slliw_T; // @[Decode.scala 49:22]
  wire  srliw = 32'h501b == _slliw_T; // @[Decode.scala 50:22]
  wire  sraiw = 32'h4000501b == _slliw_T; // @[Decode.scala 51:22]
  wire  jalr = 32'h67 == _addi_T; // @[Decode.scala 52:22]
  wire  lb = 32'h3 == _addi_T; // @[Decode.scala 53:22]
  wire  lh = 32'h1003 == _addi_T; // @[Decode.scala 54:22]
  wire  lw = 32'h2003 == _addi_T; // @[Decode.scala 55:22]
  wire  ld = 32'h3003 == _addi_T; // @[Decode.scala 56:22]
  wire  lbu = 32'h4003 == _addi_T; // @[Decode.scala 57:22]
  wire  lhu = 32'h5003 == _addi_T; // @[Decode.scala 58:22]
  wire  lwu = 32'h6003 == _addi_T; // @[Decode.scala 59:22]
  wire  csrrw = 32'h1073 == _addi_T; // @[Decode.scala 60:22]
  wire  csrrs = 32'h2073 == _addi_T; // @[Decode.scala 61:22]
  wire  ecall = 32'h73 == io_in_inst; // @[Decode.scala 62:22]
  wire  csrrc = 32'h3073 == _addi_T; // @[Decode.scala 63:22]
  wire  csrrsi = 32'h6073 == _addi_T; // @[Decode.scala 64:22]
  wire  csrrci = 32'h7073 == _addi_T; // @[Decode.scala 65:22]
  wire  _typeI_T_5 = addi | andi | xori | ori | slli | srli | srai; // @[Decode.scala 66:71]
  wire  _typeI_T_11 = _typeI_T_5 | slti | sltiu | addiw | slliw | srliw | sraiw; // @[Decode.scala 67:71]
  wire  _typeI_T_17 = _typeI_T_11 | lb | lh | lw | ld | lbu | lhu; // @[Decode.scala 68:71]
  wire  _typeI_T_23 = _typeI_T_17 | lwu | csrrw | csrrs | ecall | csrrc | csrrsi; // @[Decode.scala 69:71]
  wire  typeI = _typeI_T_23 | csrrci; // @[Decode.scala 70:24]
  wire [31:0] _auipc_T = io_in_inst & 32'h7f; // @[Decode.scala 72:22]
  wire  auipc = 32'h17 == _auipc_T; // @[Decode.scala 72:22]
  wire  lui = 32'h37 == _auipc_T; // @[Decode.scala 73:22]
  wire  typeU = auipc | lui; // @[Decode.scala 74:22]
  wire  jal = 32'h6f == _auipc_T; // @[Decode.scala 76:22]
  wire  typeJ = jal | jalr; // @[Decode.scala 77:21]
  wire  add = 32'h33 == _slliw_T; // @[Decode.scala 79:22]
  wire  sub = 32'h40000033 == _slliw_T; // @[Decode.scala 80:22]
  wire  sll = 32'h1033 == _slliw_T; // @[Decode.scala 81:22]
  wire  slt = 32'h2033 == _slliw_T; // @[Decode.scala 82:22]
  wire  sltu = 32'h3033 == _slliw_T; // @[Decode.scala 83:22]
  wire  xor_ = 32'h4033 == _slliw_T; // @[Decode.scala 84:22]
  wire  srl = 32'h5033 == _slliw_T; // @[Decode.scala 85:22]
  wire  sra = 32'h40005033 == _slliw_T; // @[Decode.scala 86:22]
  wire  or_ = 32'h6033 == _slliw_T; // @[Decode.scala 87:22]
  wire  and_ = 32'h7033 == _slliw_T; // @[Decode.scala 88:22]
  wire  addw = 32'h3b == _slliw_T; // @[Decode.scala 89:22]
  wire  subw = 32'h4000003b == _slliw_T; // @[Decode.scala 90:22]
  wire  sllw = 32'h103b == _slliw_T; // @[Decode.scala 91:22]
  wire  srlw = 32'h503b == _slliw_T; // @[Decode.scala 92:22]
  wire  sraw = 32'h4000503b == _slliw_T; // @[Decode.scala 93:22]
  wire  mret = 32'h30200073 == io_in_inst; // @[Decode.scala 94:22]
  wire  _typeR_T_4 = add | sub | sll | slt | sltu | xor_; // @[Decode.scala 95:54]
  wire  _typeR_T_9 = _typeR_T_4 | srl | sra | or_ | and_ | addw; // @[Decode.scala 96:54]
  wire  typeR = _typeR_T_9 | subw | sllw | srlw | sraw | mret; // @[Decode.scala 97:54]
  wire  beq = 32'h63 == _addi_T; // @[Decode.scala 100:22]
  wire  bne = 32'h1063 == _addi_T; // @[Decode.scala 101:22]
  wire  blt = 32'h4063 == _addi_T; // @[Decode.scala 102:22]
  wire  bge = 32'h5063 == _addi_T; // @[Decode.scala 103:22]
  wire  bltu = 32'h6063 == _addi_T; // @[Decode.scala 104:22]
  wire  bgeu = 32'h7063 == _addi_T; // @[Decode.scala 105:22]
  wire  _typeB_T_2 = beq | bne | blt | bge; // @[Decode.scala 106:38]
  wire  typeB = _typeB_T_2 | bltu | bgeu; // @[Decode.scala 107:30]
  wire  sb = 32'h23 == _addi_T; // @[Decode.scala 109:22]
  wire  sh = 32'h1023 == _addi_T; // @[Decode.scala 110:22]
  wire  sw = 32'h2023 == _addi_T; // @[Decode.scala 111:22]
  wire  sd = 32'h3023 == _addi_T; // @[Decode.scala 112:22]
  wire  _typeS_T_1 = sb | sh | sw; // @[Decode.scala 113:26]
  wire  typeS = _typeS_T_1 | sd; // @[Decode.scala 114:20]
  wire  my_inst = 32'h7b == io_in_inst; // @[Decode.scala 116:22]
  wire [51:0] imm_i_hi = io_in_inst[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [11:0] imm_i_lo = io_in_inst[31:20]; // @[Decode.scala 118:43]
  wire [63:0] imm_i = {imm_i_hi,imm_i_lo}; // @[Cat.scala 30:58]
  wire [31:0] imm_u_hi_hi = io_in_inst[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [19:0] imm_u_hi_lo = io_in_inst[31:12]; // @[Decode.scala 119:43]
  wire [63:0] imm_u = {imm_u_hi_hi,imm_u_hi_lo,12'h0}; // @[Cat.scala 30:58]
  wire [42:0] imm_j_hi_hi_hi = io_in_inst[31] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 72:12]
  wire [7:0] imm_j_hi_lo = io_in_inst[19:12]; // @[Decode.scala 120:53]
  wire  imm_j_lo_hi_hi = io_in_inst[20]; // @[Decode.scala 120:67]
  wire [9:0] imm_j_lo_hi_lo = io_in_inst[30:21]; // @[Decode.scala 120:77]
  wire [63:0] imm_j = {imm_j_hi_hi_hi,io_in_inst[31],imm_j_hi_lo,imm_j_lo_hi_hi,imm_j_lo_hi_lo,1'h0}; // @[Cat.scala 30:58]
  wire  imm_b_hi_lo = io_in_inst[7]; // @[Decode.scala 121:53]
  wire [5:0] imm_b_lo_hi_hi = io_in_inst[30:25]; // @[Decode.scala 121:62]
  wire [3:0] imm_b_lo_hi_lo = io_in_inst[11:8]; // @[Decode.scala 121:76]
  wire [55:0] imm_b = {imm_j_hi_hi_hi,io_in_inst[31],imm_b_hi_lo,imm_b_lo_hi_hi,imm_b_lo_hi_lo,1'h0}; // @[Cat.scala 30:58]
  wire [6:0] imm_s_hi_lo = io_in_inst[31:25]; // @[Decode.scala 122:43]
  wire [4:0] imm_s_lo = io_in_inst[11:7]; // @[Decode.scala 122:57]
  wire [63:0] imm_s = {imm_i_hi,imm_s_hi_lo,imm_s_lo}; // @[Cat.scala 30:58]
  wire  _alu_add_T_4 = addi | addiw | jalr | lb | lbu | lh; // @[Decode.scala 124:57]
  wire  _alu_add_T_9 = _alu_add_T_4 | lhu | lw | lwu | ld | sb; // @[Decode.scala 125:57]
  wire  _alu_add_T_14 = _alu_add_T_9 | sh | sw | sd | auipc | lui; // @[Decode.scala 126:57]
  wire  alu_add = _alu_add_T_14 | jal | add | addw; // @[Decode.scala 127:41]
  wire  alu_and = andi | and_; // @[Decode.scala 128:24]
  wire  alu_sub = subw | sub; // @[Decode.scala 129:24]
  wire  alu_slt = slti | slt; // @[Decode.scala 130:24]
  wire  alu_sltu = sltu | sltiu; // @[Decode.scala 131:24]
  wire  alu_xor = xori | xor_; // @[Decode.scala 132:24]
  wire  alu_or = ori | or_; // @[Decode.scala 133:24]
  wire  alu_sll = slli | slliw | sll | sllw; // @[Decode.scala 134:40]
  wire  alu_srl = srli | srliw | srl | srlw; // @[Decode.scala 135:40]
  wire  alu_sra = srai | sraiw | sra | sraw; // @[Decode.scala 136:40]
  wire [4:0] rs1_addr = my_inst ? 5'ha : io_in_inst[19:15]; // @[Decode.scala 138:22]
  wire [4:0] rs2_addr = io_in_inst[24:20]; // @[Decode.scala 139:23]
  wire  rs1_en = ~(ecall | auipc | lui | jal); // @[Decode.scala 140:19]
  wire  rs2_en = typeR | typeB | typeS; // @[Decode.scala 141:34]
  wire  t_int = io_time_int & io_in_valid; // @[Decode.scala 150:33]
  wire  _rs1_forward_T_1 = rs1_addr == io_ex_wdest; // @[Decode.scala 152:53]
  wire  rs1_forward = rs1_addr != 5'h0 & (rs1_addr == io_ex_wdest | rs1_addr == io_wb_wdest) & rs1_en; // @[Decode.scala 152:92]
  wire  _rs2_forward_T_1 = rs2_addr == io_ex_wdest; // @[Decode.scala 153:53]
  wire  rs2_forward = rs2_addr != 5'h0 & (rs2_addr == io_ex_wdest | rs2_addr == io_wb_wdest) & rs2_en; // @[Decode.scala 153:92]
  wire [63:0] _rs1_value_T_1 = _rs1_forward_T_1 ? io_ex_result : io_wb_result; // @[Decode.scala 154:41]
  wire [63:0] rs1_value = rs1_forward ? _rs1_value_T_1 : io_rs1_data; // @[Decode.scala 154:24]
  wire [63:0] _rs2_value_T_1 = _rs2_forward_T_1 ? io_ex_result : io_wb_result; // @[Decode.scala 155:41]
  wire [63:0] rs2_value = rs2_forward ? _rs2_value_T_1 : io_rs2_data; // @[Decode.scala 155:24]
  wire  id_wen = ~(ecall | mret | my_inst | typeS | typeB); // @[Decode.scala 157:19]
  wire [5:0] _id_opcode_T_1 = typeI ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [5:0] _id_opcode_T_2 = _id_opcode_T_1 & 6'h10; // @[Decode.scala 160:47]
  wire [5:0] _id_opcode_T_4 = typeU ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [5:0] _id_opcode_T_5 = _id_opcode_T_4 & 6'h20; // @[Decode.scala 161:47]
  wire [5:0] _id_opcode_T_6 = _id_opcode_T_2 | _id_opcode_T_5; // @[Decode.scala 160:64]
  wire [5:0] _id_opcode_T_8 = typeJ ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [5:0] _id_opcode_T_9 = _id_opcode_T_8 & 6'h2; // @[Decode.scala 162:47]
  wire [5:0] _id_opcode_T_10 = _id_opcode_T_6 | _id_opcode_T_9; // @[Decode.scala 161:64]
  wire [5:0] _id_opcode_T_12 = typeR ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [5:0] _id_opcode_T_13 = _id_opcode_T_12 & 6'h8; // @[Decode.scala 163:47]
  wire [5:0] _id_opcode_T_14 = _id_opcode_T_10 | _id_opcode_T_13; // @[Decode.scala 162:64]
  wire [5:0] _id_opcode_T_16 = typeB ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [5:0] _id_opcode_T_17 = _id_opcode_T_16 & 6'h1; // @[Decode.scala 164:47]
  wire [5:0] _id_opcode_T_18 = _id_opcode_T_14 | _id_opcode_T_17; // @[Decode.scala 163:64]
  wire [5:0] _id_opcode_T_20 = typeS ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [5:0] _id_opcode_T_21 = _id_opcode_T_20 & 6'h4; // @[Decode.scala 165:47]
  wire [5:0] id_opcode = _id_opcode_T_18 | _id_opcode_T_21; // @[Decode.scala 164:64]
  wire [11:0] _id_aluop_T_1 = alu_add ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _id_aluop_T_2 = _id_aluop_T_1 & 12'h1; // @[Decode.scala 166:49]
  wire [11:0] _id_aluop_T_4 = alu_and ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _id_aluop_T_5 = _id_aluop_T_4 & 12'h40; // @[Decode.scala 167:49]
  wire [11:0] _id_aluop_T_6 = _id_aluop_T_2 | _id_aluop_T_5; // @[Decode.scala 166:68]
  wire [11:0] _id_aluop_T_8 = alu_or ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _id_aluop_T_9 = _id_aluop_T_8 & 12'h20; // @[Decode.scala 168:49]
  wire [11:0] _id_aluop_T_10 = _id_aluop_T_6 | _id_aluop_T_9; // @[Decode.scala 167:68]
  wire [11:0] _id_aluop_T_12 = alu_sll ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _id_aluop_T_13 = _id_aluop_T_12 & 12'h80; // @[Decode.scala 169:49]
  wire [11:0] _id_aluop_T_14 = _id_aluop_T_10 | _id_aluop_T_13; // @[Decode.scala 168:68]
  wire [11:0] _id_aluop_T_16 = alu_slt ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _id_aluop_T_17 = _id_aluop_T_16 & 12'h4; // @[Decode.scala 170:49]
  wire [11:0] _id_aluop_T_18 = _id_aluop_T_14 | _id_aluop_T_17; // @[Decode.scala 169:68]
  wire [11:0] _id_aluop_T_20 = alu_sltu ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _id_aluop_T_21 = _id_aluop_T_20 & 12'h8; // @[Decode.scala 171:49]
  wire [11:0] _id_aluop_T_22 = _id_aluop_T_18 | _id_aluop_T_21; // @[Decode.scala 170:68]
  wire [11:0] _id_aluop_T_24 = alu_sra ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _id_aluop_T_25 = _id_aluop_T_24 & 12'h200; // @[Decode.scala 172:49]
  wire [11:0] _id_aluop_T_26 = _id_aluop_T_22 | _id_aluop_T_25; // @[Decode.scala 171:68]
  wire [11:0] _id_aluop_T_28 = alu_srl ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _id_aluop_T_29 = _id_aluop_T_28 & 12'h100; // @[Decode.scala 173:49]
  wire [11:0] _id_aluop_T_30 = _id_aluop_T_26 | _id_aluop_T_29; // @[Decode.scala 172:68]
  wire [11:0] _id_aluop_T_32 = alu_sub ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _id_aluop_T_33 = _id_aluop_T_32 & 12'h2; // @[Decode.scala 174:49]
  wire [11:0] _id_aluop_T_34 = _id_aluop_T_30 | _id_aluop_T_33; // @[Decode.scala 173:68]
  wire [11:0] _id_aluop_T_36 = alu_xor ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _id_aluop_T_37 = _id_aluop_T_36 & 12'h10; // @[Decode.scala 175:49]
  wire [6:0] _id_loadop_T_1 = lb ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [6:0] _id_loadop_T_2 = _id_loadop_T_1 & 7'h1; // @[Decode.scala 176:45]
  wire [6:0] _id_loadop_T_4 = lh ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [6:0] _id_loadop_T_5 = _id_loadop_T_4 & 7'h4; // @[Decode.scala 177:45]
  wire [6:0] _id_loadop_T_6 = _id_loadop_T_2 | _id_loadop_T_5; // @[Decode.scala 176:64]
  wire [6:0] _id_loadop_T_8 = lw ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [6:0] _id_loadop_T_9 = _id_loadop_T_8 & 7'h10; // @[Decode.scala 178:45]
  wire [6:0] _id_loadop_T_10 = _id_loadop_T_6 | _id_loadop_T_9; // @[Decode.scala 177:64]
  wire [6:0] _id_loadop_T_12 = ld ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [6:0] _id_loadop_T_13 = _id_loadop_T_12 & 7'h40; // @[Decode.scala 179:45]
  wire [6:0] _id_loadop_T_14 = _id_loadop_T_10 | _id_loadop_T_13; // @[Decode.scala 178:64]
  wire [6:0] _id_loadop_T_16 = lbu ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [6:0] _id_loadop_T_17 = _id_loadop_T_16 & 7'h2; // @[Decode.scala 180:45]
  wire [6:0] _id_loadop_T_18 = _id_loadop_T_14 | _id_loadop_T_17; // @[Decode.scala 179:64]
  wire [6:0] _id_loadop_T_20 = lhu ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [6:0] _id_loadop_T_21 = _id_loadop_T_20 & 7'h8; // @[Decode.scala 181:45]
  wire [6:0] _id_loadop_T_22 = _id_loadop_T_18 | _id_loadop_T_21; // @[Decode.scala 180:64]
  wire [6:0] _id_loadop_T_24 = lwu ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [6:0] _id_loadop_T_25 = _id_loadop_T_24 & 7'h20; // @[Decode.scala 182:45]
  wire [3:0] _id_storeop_T_1 = sb ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _id_storeop_T_2 = _id_storeop_T_1 & 4'h1; // @[Decode.scala 183:45]
  wire [3:0] _id_storeop_T_4 = sh ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _id_storeop_T_5 = _id_storeop_T_4 & 4'h2; // @[Decode.scala 184:45]
  wire [3:0] _id_storeop_T_6 = _id_storeop_T_2 | _id_storeop_T_5; // @[Decode.scala 183:64]
  wire [3:0] _id_storeop_T_8 = sw ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _id_storeop_T_9 = _id_storeop_T_8 & 4'h4; // @[Decode.scala 185:45]
  wire [3:0] _id_storeop_T_10 = _id_storeop_T_6 | _id_storeop_T_9; // @[Decode.scala 184:64]
  wire [3:0] _id_storeop_T_12 = sd ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _id_storeop_T_13 = _id_storeop_T_12 & 4'h8; // @[Decode.scala 186:45]
  wire [3:0] _id_sysop_T_1 = csrrs ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _id_sysop_T_2 = _id_sysop_T_1 & 4'h2; // @[Decode.scala 187:47]
  wire [3:0] _id_sysop_T_4 = csrrsi ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _id_sysop_T_5 = _id_sysop_T_4 & 4'h8; // @[Decode.scala 188:47]
  wire [3:0] _id_sysop_T_6 = _id_sysop_T_2 | _id_sysop_T_5; // @[Decode.scala 187:68]
  wire [3:0] _id_sysop_T_8 = csrrc ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _id_sysop_T_9 = _id_sysop_T_8 & 4'h3; // @[Decode.scala 189:47]
  wire [3:0] _id_sysop_T_10 = _id_sysop_T_6 | _id_sysop_T_9; // @[Decode.scala 188:68]
  wire [3:0] _id_sysop_T_12 = csrrci ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _id_sysop_T_13 = _id_sysop_T_12 & 4'h9; // @[Decode.scala 190:47]
  wire [3:0] _id_sysop_T_14 = _id_sysop_T_10 | _id_sysop_T_13; // @[Decode.scala 189:68]
  wire [3:0] _id_sysop_T_16 = csrrw ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _id_sysop_T_17 = _id_sysop_T_16 & 4'h1; // @[Decode.scala 191:47]
  wire [3:0] _id_sysop_T_18 = _id_sysop_T_14 | _id_sysop_T_17; // @[Decode.scala 190:68]
  wire [3:0] _id_sysop_T_20 = ecall ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _id_sysop_T_21 = _id_sysop_T_20 & 4'h4; // @[Decode.scala 192:47]
  wire [3:0] _id_sysop_T_22 = _id_sysop_T_18 | _id_sysop_T_21; // @[Decode.scala 191:68]
  wire [3:0] _id_sysop_T_24 = mret ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _id_sysop_T_25 = _id_sysop_T_24 & 4'h5; // @[Decode.scala 193:47]
  wire [3:0] _id_sysop_T_26 = _id_sysop_T_22 | _id_sysop_T_25; // @[Decode.scala 192:68]
  wire [3:0] _id_sysop_T_28 = t_int ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _id_sysop_T_29 = _id_sysop_T_28 & 4'h7; // @[Decode.scala 194:47]
  wire [31:0] _id_op1_T_2 = auipc ? io_in_pc : 32'h0; // @[Decode.scala 197:41]
  wire [63:0] _id_op1_T_4 = 6'h10 == id_opcode ? rs1_value : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _id_op1_T_6 = 6'h20 == id_opcode ? {{32'd0}, _id_op1_T_2} : _id_op1_T_4; // @[Mux.scala 80:57]
  wire [63:0] _id_op1_T_8 = 6'h2 == id_opcode ? {{32'd0}, io_in_pc} : _id_op1_T_6; // @[Mux.scala 80:57]
  wire [63:0] _id_op1_T_10 = 6'h8 == id_opcode ? rs1_value : _id_op1_T_8; // @[Mux.scala 80:57]
  wire [63:0] _id_op1_T_12 = 6'h1 == id_opcode ? rs1_value : _id_op1_T_10; // @[Mux.scala 80:57]
  wire [63:0] id_op1 = 6'h4 == id_opcode ? rs1_value : _id_op1_T_12; // @[Mux.scala 80:57]
  wire [63:0] _id_op2_T_1 = 6'h10 == id_opcode ? imm_i : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _id_op2_T_3 = 6'h20 == id_opcode ? imm_u : _id_op2_T_1; // @[Mux.scala 80:57]
  wire [63:0] _id_op2_T_5 = 6'h2 == id_opcode ? 64'h4 : _id_op2_T_3; // @[Mux.scala 80:57]
  wire [63:0] _id_op2_T_7 = 6'h8 == id_opcode ? rs2_value : _id_op2_T_5; // @[Mux.scala 80:57]
  wire [63:0] _id_op2_T_9 = 6'h1 == id_opcode ? rs2_value : _id_op2_T_7; // @[Mux.scala 80:57]
  wire  _id_typew_T_4 = addiw | slliw | srliw | sraiw | addw | subw; // @[Decode.scala 211:60]
  wire [10:0] _redirectop_T_1 = jal ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _redirectop_T_2 = _redirectop_T_1 & 11'h10; // @[Decode.scala 218:52]
  wire [10:0] _redirectop_T_4 = jalr ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _redirectop_T_5 = _redirectop_T_4 & 11'h8; // @[Decode.scala 219:52]
  wire [10:0] _redirectop_T_6 = _redirectop_T_2 | _redirectop_T_5; // @[Decode.scala 218:77]
  wire [10:0] _redirectop_T_8 = beq ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _redirectop_T_9 = _redirectop_T_8 & 11'h400; // @[Decode.scala 220:52]
  wire [10:0] _redirectop_T_10 = _redirectop_T_6 | _redirectop_T_9; // @[Decode.scala 219:77]
  wire [10:0] _redirectop_T_12 = bne ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _redirectop_T_13 = _redirectop_T_12 & 11'h200; // @[Decode.scala 221:52]
  wire [10:0] _redirectop_T_14 = _redirectop_T_10 | _redirectop_T_13; // @[Decode.scala 220:77]
  wire [10:0] _redirectop_T_16 = blt ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _redirectop_T_17 = _redirectop_T_16 & 11'h100; // @[Decode.scala 222:52]
  wire [10:0] _redirectop_T_18 = _redirectop_T_14 | _redirectop_T_17; // @[Decode.scala 221:77]
  wire [10:0] _redirectop_T_20 = bge ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _redirectop_T_21 = _redirectop_T_20 & 11'h80; // @[Decode.scala 223:52]
  wire [10:0] _redirectop_T_22 = _redirectop_T_18 | _redirectop_T_21; // @[Decode.scala 222:77]
  wire [10:0] _redirectop_T_24 = bltu ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _redirectop_T_25 = _redirectop_T_24 & 11'h40; // @[Decode.scala 224:52]
  wire [10:0] _redirectop_T_26 = _redirectop_T_22 | _redirectop_T_25; // @[Decode.scala 223:77]
  wire [10:0] _redirectop_T_28 = bgeu ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _redirectop_T_29 = _redirectop_T_28 & 11'h20; // @[Decode.scala 225:52]
  wire [10:0] _redirectop_T_30 = _redirectop_T_26 | _redirectop_T_29; // @[Decode.scala 224:77]
  wire [10:0] _redirectop_T_32 = ecall ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _redirectop_T_33 = _redirectop_T_32 & 11'h4; // @[Decode.scala 226:52]
  wire [10:0] _redirectop_T_34 = _redirectop_T_30 | _redirectop_T_33; // @[Decode.scala 225:77]
  wire [10:0] _redirectop_T_36 = mret ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _redirectop_T_37 = _redirectop_T_36 & 11'h2; // @[Decode.scala 227:52]
  wire [10:0] _redirectop_T_38 = _redirectop_T_34 | _redirectop_T_37; // @[Decode.scala 226:77]
  wire [10:0] _redirectop_T_40 = t_int ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _redirectop_T_41 = _redirectop_T_40 & 11'h1; // @[Decode.scala 228:52]
  wire [10:0] redirectop = _redirectop_T_38 | _redirectop_T_41; // @[Decode.scala 227:77]
  wire  br_stall = io_stall & (rs1_forward | rs2_forward); // @[Decode.scala 239:30]
  wire [63:0] _GEN_0 = {{32'd0}, io_in_bp_targer}; // @[Decode.scala 243:60]
  wire  _mis_predict_T_4 = ctrl_io_jmp ? io_in_bp_taken & ctrl_io_target != _GEN_0 | ~io_in_bp_taken : io_in_bp_taken; // @[Decode.scala 243:24]
  wire  mis_predict = _mis_predict_T_4 & ~br_stall; // @[Decode.scala 243:109]
  Ctrl ctrl ( // @[Decode.scala 217:20]
    .io_redirectop(ctrl_io_redirectop),
    .io_pc(ctrl_io_pc),
    .io_imm_i(ctrl_io_imm_i),
    .io_imm_j(ctrl_io_imm_j),
    .io_imm_b(ctrl_io_imm_b),
    .io_rs1_value(ctrl_io_rs1_value),
    .io_rs2_value(ctrl_io_rs2_value),
    .io_mtvec(ctrl_io_mtvec),
    .io_mepc(ctrl_io_mepc),
    .io_jmp(ctrl_io_jmp),
    .io_target(ctrl_io_target)
  );
  assign io_rs1_addr = my_inst ? 5'ha : io_in_inst[19:15]; // @[Decode.scala 138:22]
  assign io_rs2_addr = io_in_inst[24:20]; // @[Decode.scala 139:23]
  assign io_out_valid = io_in_valid; // @[Decode.scala 255:21]
  assign io_out_pc = io_in_pc; // @[Decode.scala 256:21]
  assign io_out_inst = io_in_inst; // @[Decode.scala 257:21]
  assign io_out_wen = ~(ecall | mret | my_inst | typeS | typeB); // @[Decode.scala 157:19]
  assign io_out_wdest = id_wen ? imm_s_lo : 5'h0; // @[Decode.scala 158:22]
  assign io_out_op1 = my_inst ? rs1_value : id_op1; // @[Decode.scala 261:27]
  assign io_out_op2 = 6'h4 == id_opcode ? imm_s : _id_op2_T_9; // @[Mux.scala 80:57]
  assign io_out_typew = _id_typew_T_4 | sllw | srlw | sraw; // @[Decode.scala 212:43]
  assign io_out_wmem = rs2_forward ? _rs2_value_T_1 : io_rs2_data; // @[Decode.scala 155:24]
  assign io_out_aluop = _id_aluop_T_34 | _id_aluop_T_37; // @[Decode.scala 174:68]
  assign io_out_loadop = _id_loadop_T_22 | _id_loadop_T_25; // @[Decode.scala 181:64]
  assign io_out_storeop = _id_storeop_T_10 | _id_storeop_T_13; // @[Decode.scala 185:64]
  assign io_out_sysop = _id_sysop_T_26 | _id_sysop_T_29; // @[Decode.scala 193:68]
  assign io_jmp_packet_valid = redirectop != 11'h0; // @[Decode.scala 245:39]
  assign io_jmp_packet_inst_pc = io_in_pc; // @[Decode.scala 246:25]
  assign io_jmp_packet_jmp = ctrl_io_jmp; // @[Decode.scala 247:25]
  assign io_jmp_packet_jmp_pc = ctrl_io_target[31:0]; // @[Decode.scala 248:25]
  assign io_jmp_packet_mis = io_jmp_packet_valid & mis_predict; // @[Decode.scala 249:48]
  assign ctrl_io_redirectop = _redirectop_T_38 | _redirectop_T_41; // @[Decode.scala 227:77]
  assign ctrl_io_pc = io_in_pc; // @[Decode.scala 230:22]
  assign ctrl_io_imm_i = imm_i[31:0]; // @[Decode.scala 231:22]
  assign ctrl_io_imm_j = imm_j[31:0]; // @[Decode.scala 232:22]
  assign ctrl_io_imm_b = imm_b[31:0]; // @[Decode.scala 233:22]
  assign ctrl_io_rs1_value = rs1_forward ? _rs1_value_T_1 : io_rs1_data; // @[Decode.scala 154:24]
  assign ctrl_io_rs2_value = rs2_forward ? _rs2_value_T_1 : io_rs2_data; // @[Decode.scala 155:24]
  assign ctrl_io_mtvec = io_mtvec; // @[Decode.scala 236:22]
  assign ctrl_io_mepc = io_mepc; // @[Decode.scala 237:22]
endmodule
module Execution(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_wen,
  input  [4:0]  io_in_wdest,
  input  [63:0] io_in_op1,
  input  [63:0] io_in_op2,
  input         io_in_typew,
  input  [63:0] io_in_wmem,
  input  [11:0] io_in_aluop,
  input  [6:0]  io_in_loadop,
  input  [3:0]  io_in_storeop,
  input  [3:0]  io_in_sysop,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_wen,
  output [4:0]  io_out_wdest,
  output [63:0] io_out_wdata,
  output [63:0] io_out_op1,
  output [63:0] io_out_op2,
  output        io_out_typew,
  output [63:0] io_out_wmem,
  output [31:0] io_out_mem_addr,
  output [11:0] io_out_aluop,
  output [6:0]  io_out_loadop,
  output [3:0]  io_out_storeop,
  output [3:0]  io_out_sysop,
  output        io_busy,
  output [11:0] io_csr_raddr,
  input  [63:0] io_csr_rdata,
  output        io_dmem_data_valid,
  input         io_dmem_data_ready,
  output        io_dmem_data_req,
  output [31:0] io_dmem_data_addr,
  output [1:0]  io_dmem_data_size,
  output [7:0]  io_dmem_data_strb,
  input  [63:0] io_dmem_data_read,
  output [63:0] io_dmem_data_write,
  output        io_cmp_ren,
  output        io_cmp_wen,
  output [63:0] io_cmp_addr,
  output [63:0] io_cmp_wdata,
  input  [63:0] io_cmp_rdata,
  output [4:0]  io_ex_wdest,
  output [63:0] io_ex_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] in1_hi = io_in_op1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] in1_lo = io_in_op1[31:0]; // @[Execution.scala 44:92]
  wire [63:0] _in1_T_3 = {in1_hi,in1_lo}; // @[Cat.scala 30:58]
  wire [63:0] _in1_T_4 = {32'h0,in1_lo}; // @[Cat.scala 30:58]
  wire [63:0] _in1_T_5 = io_in_aluop == 12'h200 ? _in1_T_3 : _in1_T_4; // @[Execution.scala 44:30]
  wire [63:0] in1 = io_in_typew ? _in1_T_5 : io_in_op1; // @[Execution.scala 44:16]
  wire [5:0] shamt = io_in_typew ? {{1'd0}, io_in_op2[4:0]} : io_in_op2[5:0]; // @[Execution.scala 47:15]
  wire [63:0] _alu_result_0_T_1 = in1 + io_in_op2; // @[Execution.scala 50:29]
  wire [63:0] _alu_result_0_T_3 = in1 - io_in_op2; // @[Execution.scala 51:29]
  wire [63:0] _alu_result_0_T_4 = io_in_typew ? _in1_T_5 : io_in_op1; // @[Execution.scala 52:35]
  wire  _alu_result_0_T_6 = $signed(_alu_result_0_T_4) < $signed(io_in_op2); // @[Execution.scala 52:38]
  wire  _alu_result_0_T_7 = in1 < io_in_op2; // @[Execution.scala 53:29]
  wire [63:0] _alu_result_0_T_8 = in1 ^ io_in_op2; // @[Execution.scala 54:29]
  wire [63:0] _alu_result_0_T_9 = in1 | io_in_op2; // @[Execution.scala 55:29]
  wire [63:0] _alu_result_0_T_10 = in1 & io_in_op2; // @[Execution.scala 56:29]
  wire [126:0] _GEN_8 = {{63'd0}, in1}; // @[Execution.scala 57:30]
  wire [126:0] _alu_result_0_T_11 = _GEN_8 << shamt; // @[Execution.scala 57:30]
  wire [63:0] _alu_result_0_T_13 = in1 >> shamt; // @[Execution.scala 58:29]
  wire [63:0] _alu_result_0_T_16 = $signed(_alu_result_0_T_4) >>> shamt; // @[Execution.scala 59:54]
  wire [63:0] _alu_result_0_T_18 = 12'h1 == io_in_aluop ? _alu_result_0_T_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_20 = 12'h2 == io_in_aluop ? _alu_result_0_T_3 : _alu_result_0_T_18; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_22 = 12'h4 == io_in_aluop ? {{63'd0}, _alu_result_0_T_6} : _alu_result_0_T_20; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_24 = 12'h8 == io_in_aluop ? {{63'd0}, _alu_result_0_T_7} : _alu_result_0_T_22; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_26 = 12'h10 == io_in_aluop ? _alu_result_0_T_8 : _alu_result_0_T_24; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_28 = 12'h20 == io_in_aluop ? _alu_result_0_T_9 : _alu_result_0_T_26; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_30 = 12'h40 == io_in_aluop ? _alu_result_0_T_10 : _alu_result_0_T_28; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_32 = 12'h80 == io_in_aluop ? _alu_result_0_T_11[63:0] : _alu_result_0_T_30; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_0_T_34 = 12'h100 == io_in_aluop ? _alu_result_0_T_13 : _alu_result_0_T_32; // @[Mux.scala 80:57]
  wire [63:0] alu_result_0 = 12'h200 == io_in_aluop ? _alu_result_0_T_16 : _alu_result_0_T_34; // @[Mux.scala 80:57]
  wire [31:0] alu_result_hi = alu_result_0[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] alu_result_lo = alu_result_0[31:0]; // @[Execution.scala 61:75]
  wire [63:0] _alu_result_T_2 = {alu_result_hi,alu_result_lo}; // @[Cat.scala 30:58]
  wire [63:0] alu_result = io_in_typew ? _alu_result_T_2 : alu_result_0; // @[Execution.scala 61:20]
  wire  _cmp_ren_T = io_in_loadop != 7'h0; // @[Execution.scala 64:29]
  wire  _cmp_ren_T_3 = io_dmem_data_addr == 32'h2004000 | io_dmem_data_addr == 32'h200bff8; // @[Execution.scala 64:79]
  wire  cmp_ren = io_in_loadop != 7'h0 & (io_dmem_data_addr == 32'h2004000 | io_dmem_data_addr == 32'h200bff8); // @[Execution.scala 64:38]
  wire  _cmp_wen_T = io_in_storeop != 4'h0; // @[Execution.scala 65:30]
  wire  cmp_wen = io_in_storeop != 4'h0 & _cmp_ren_T_3; // @[Execution.scala 65:38]
  wire  _data_valid_T_2 = ~cmp_wen; // @[Execution.scala 80:59]
  wire  data_valid = (_cmp_ren_T | _cmp_wen_T) & (~cmp_ren & ~cmp_wen); // @[Execution.scala 80:43]
  wire [63:0] data_read = cmp_ren ? io_cmp_rdata : io_dmem_data_read; // @[Execution.scala 83:24]
  wire [55:0] mem_wdata_lb_hi = data_read[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mem_wdata_lb_lo = data_read[7:0]; // @[Execution.scala 86:60]
  wire [63:0] mem_wdata_lb = {mem_wdata_lb_hi,mem_wdata_lb_lo}; // @[Cat.scala 30:58]
  wire [47:0] mem_wdata_lh_hi = data_read[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [15:0] mem_wdata_lh_lo = data_read[15:0]; // @[Execution.scala 87:60]
  wire [63:0] mem_wdata_lh = {mem_wdata_lh_hi,mem_wdata_lh_lo}; // @[Cat.scala 30:58]
  wire [31:0] mem_wdata_lw_hi = data_read[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] mem_wdata_lw_lo = data_read[31:0]; // @[Execution.scala 88:60]
  wire [63:0] mem_wdata_lw = {mem_wdata_lw_hi,mem_wdata_lw_lo}; // @[Cat.scala 30:58]
  wire [63:0] mem_wdata_lbu = {56'h0,mem_wdata_lb_lo}; // @[Cat.scala 30:58]
  wire [63:0] mem_wdata_lhu = {48'h0,mem_wdata_lh_lo}; // @[Cat.scala 30:58]
  wire [63:0] mem_wdata_lwu = {32'h0,mem_wdata_lw_lo}; // @[Cat.scala 30:58]
  wire [31:0] _mem_wdata_T = io_in_inst & 32'h707f; // @[Execution.scala 93:41]
  wire  _mem_wdata_T_1 = 32'h3 == _mem_wdata_T; // @[Execution.scala 93:41]
  wire [63:0] _mem_wdata_T_3 = _mem_wdata_T_1 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_4 = _mem_wdata_T_3 & mem_wdata_lb; // @[Execution.scala 93:50]
  wire  _mem_wdata_T_6 = 32'h1003 == _mem_wdata_T; // @[Execution.scala 94:41]
  wire [63:0] _mem_wdata_T_8 = _mem_wdata_T_6 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_9 = _mem_wdata_T_8 & mem_wdata_lh; // @[Execution.scala 94:50]
  wire [63:0] _mem_wdata_T_10 = _mem_wdata_T_4 | _mem_wdata_T_9; // @[Execution.scala 93:67]
  wire  _mem_wdata_T_12 = 32'h2003 == _mem_wdata_T; // @[Execution.scala 95:41]
  wire [63:0] _mem_wdata_T_14 = _mem_wdata_T_12 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_15 = _mem_wdata_T_14 & mem_wdata_lw; // @[Execution.scala 95:50]
  wire [63:0] _mem_wdata_T_16 = _mem_wdata_T_10 | _mem_wdata_T_15; // @[Execution.scala 94:67]
  wire  _mem_wdata_T_18 = 32'h3003 == _mem_wdata_T; // @[Execution.scala 96:41]
  wire [63:0] _mem_wdata_T_20 = _mem_wdata_T_18 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_21 = _mem_wdata_T_20 & data_read; // @[Execution.scala 96:50]
  wire [63:0] _mem_wdata_T_22 = _mem_wdata_T_16 | _mem_wdata_T_21; // @[Execution.scala 95:67]
  wire  _mem_wdata_T_24 = 32'h4003 == _mem_wdata_T; // @[Execution.scala 97:41]
  wire [63:0] _mem_wdata_T_26 = _mem_wdata_T_24 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_27 = _mem_wdata_T_26 & mem_wdata_lbu; // @[Execution.scala 97:50]
  wire [63:0] _mem_wdata_T_28 = _mem_wdata_T_22 | _mem_wdata_T_27; // @[Execution.scala 96:67]
  wire  _mem_wdata_T_30 = 32'h5003 == _mem_wdata_T; // @[Execution.scala 98:41]
  wire [63:0] _mem_wdata_T_32 = _mem_wdata_T_30 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_33 = _mem_wdata_T_32 & mem_wdata_lhu; // @[Execution.scala 98:50]
  wire [63:0] _mem_wdata_T_34 = _mem_wdata_T_28 | _mem_wdata_T_33; // @[Execution.scala 97:67]
  wire  _mem_wdata_T_36 = 32'h6003 == _mem_wdata_T; // @[Execution.scala 99:41]
  wire [63:0] _mem_wdata_T_38 = _mem_wdata_T_36 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _mem_wdata_T_39 = _mem_wdata_T_38 & mem_wdata_lwu; // @[Execution.scala 99:50]
  wire [63:0] mem_wdata = _mem_wdata_T_34 | _mem_wdata_T_39; // @[Execution.scala 98:67]
  wire [7:0] data_write_sb_lo = io_in_wmem[7:0]; // @[Execution.scala 103:43]
  wire [63:0] _data_write_sb_T_1 = {56'h0,data_write_sb_lo}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_2 = {48'h0,data_write_sb_lo,8'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_3 = {40'h0,data_write_sb_lo,16'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_4 = {32'h0,data_write_sb_lo,24'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_5 = {24'h0,data_write_sb_lo,32'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_6 = {16'h0,data_write_sb_lo,40'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_7 = {8'h0,data_write_sb_lo,48'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_8 = {data_write_sb_lo,56'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sb_T_10 = 3'h1 == alu_result[2:0] ? _data_write_sb_T_2 : _data_write_sb_T_1; // @[Mux.scala 80:57]
  wire [63:0] _data_write_sb_T_12 = 3'h2 == alu_result[2:0] ? _data_write_sb_T_3 : _data_write_sb_T_10; // @[Mux.scala 80:57]
  wire [63:0] _data_write_sb_T_14 = 3'h3 == alu_result[2:0] ? _data_write_sb_T_4 : _data_write_sb_T_12; // @[Mux.scala 80:57]
  wire [63:0] _data_write_sb_T_16 = 3'h4 == alu_result[2:0] ? _data_write_sb_T_5 : _data_write_sb_T_14; // @[Mux.scala 80:57]
  wire [63:0] _data_write_sb_T_18 = 3'h5 == alu_result[2:0] ? _data_write_sb_T_6 : _data_write_sb_T_16; // @[Mux.scala 80:57]
  wire [63:0] _data_write_sb_T_20 = 3'h6 == alu_result[2:0] ? _data_write_sb_T_7 : _data_write_sb_T_18; // @[Mux.scala 80:57]
  wire [63:0] data_write_sb = 3'h7 == alu_result[2:0] ? _data_write_sb_T_8 : _data_write_sb_T_20; // @[Mux.scala 80:57]
  wire [1:0] _data_strb_sb_T_2 = 3'h1 == alu_result[2:0] ? 2'h2 : 2'h1; // @[Mux.scala 80:57]
  wire [2:0] _data_strb_sb_T_4 = 3'h2 == alu_result[2:0] ? 3'h4 : {{1'd0}, _data_strb_sb_T_2}; // @[Mux.scala 80:57]
  wire [3:0] _data_strb_sb_T_6 = 3'h3 == alu_result[2:0] ? 4'h8 : {{1'd0}, _data_strb_sb_T_4}; // @[Mux.scala 80:57]
  wire [4:0] _data_strb_sb_T_8 = 3'h4 == alu_result[2:0] ? 5'h10 : {{1'd0}, _data_strb_sb_T_6}; // @[Mux.scala 80:57]
  wire [5:0] _data_strb_sb_T_10 = 3'h5 == alu_result[2:0] ? 6'h20 : {{1'd0}, _data_strb_sb_T_8}; // @[Mux.scala 80:57]
  wire [6:0] _data_strb_sb_T_12 = 3'h6 == alu_result[2:0] ? 7'h40 : {{1'd0}, _data_strb_sb_T_10}; // @[Mux.scala 80:57]
  wire [7:0] data_strb_sb = 3'h7 == alu_result[2:0] ? 8'h80 : {{1'd0}, _data_strb_sb_T_12}; // @[Mux.scala 80:57]
  wire [15:0] data_write_sh_lo = io_in_wmem[15:0]; // @[Execution.scala 124:42]
  wire [63:0] _data_write_sh_T_1 = {48'h0,data_write_sh_lo}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sh_T_2 = {32'h0,data_write_sh_lo,16'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sh_T_3 = {16'h0,data_write_sh_lo,32'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sh_T_4 = {data_write_sh_lo,48'h0}; // @[Cat.scala 30:58]
  wire [63:0] _data_write_sh_T_6 = 2'h1 == alu_result[2:1] ? _data_write_sh_T_2 : _data_write_sh_T_1; // @[Mux.scala 80:57]
  wire [63:0] _data_write_sh_T_8 = 2'h2 == alu_result[2:1] ? _data_write_sh_T_3 : _data_write_sh_T_6; // @[Mux.scala 80:57]
  wire [63:0] data_write_sh = 2'h3 == alu_result[2:1] ? _data_write_sh_T_4 : _data_write_sh_T_8; // @[Mux.scala 80:57]
  wire [3:0] _data_strb_sh_T_2 = 2'h1 == alu_result[2:1] ? 4'hc : 4'h3; // @[Mux.scala 80:57]
  wire [5:0] _data_strb_sh_T_4 = 2'h2 == alu_result[2:1] ? 6'h30 : {{2'd0}, _data_strb_sh_T_2}; // @[Mux.scala 80:57]
  wire [7:0] data_strb_sh = 2'h3 == alu_result[2:1] ? 8'hc0 : {{2'd0}, _data_strb_sh_T_4}; // @[Mux.scala 80:57]
  wire [32:0] data_write_sw_lo = io_in_wmem[32:0]; // @[Execution.scala 137:41]
  wire [64:0] _data_write_sw_T_1 = {32'h0,data_write_sw_lo}; // @[Cat.scala 30:58]
  wire [64:0] _data_write_sw_T_2 = {data_write_sw_lo,32'h0}; // @[Cat.scala 30:58]
  wire [64:0] data_write_sw = alu_result[2] ? _data_write_sw_T_2 : _data_write_sw_T_1; // @[Mux.scala 80:57]
  wire [7:0] data_strb_sw = alu_result[2] ? 8'hf0 : 8'hf; // @[Mux.scala 80:57]
  wire  _data_write_T_1 = 32'h3023 == _mem_wdata_T; // @[Execution.scala 147:39]
  wire [63:0] _data_write_T_3 = _data_write_T_1 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _data_write_T_4 = _data_write_T_3 & io_in_wmem; // @[Execution.scala 147:47]
  wire  _data_write_T_6 = 32'h2023 == _mem_wdata_T; // @[Execution.scala 148:39]
  wire [63:0] _data_write_T_8 = _data_write_T_6 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [64:0] _GEN_9 = {{1'd0}, _data_write_T_8}; // @[Execution.scala 148:47]
  wire [64:0] _data_write_T_9 = _GEN_9 & data_write_sw; // @[Execution.scala 148:47]
  wire [64:0] _GEN_10 = {{1'd0}, _data_write_T_4}; // @[Execution.scala 147:64]
  wire [64:0] _data_write_T_10 = _GEN_10 | _data_write_T_9; // @[Execution.scala 147:64]
  wire  _data_write_T_12 = 32'h1023 == _mem_wdata_T; // @[Execution.scala 149:39]
  wire [63:0] _data_write_T_14 = _data_write_T_12 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _data_write_T_15 = _data_write_T_14 & data_write_sh; // @[Execution.scala 149:47]
  wire [64:0] _GEN_11 = {{1'd0}, _data_write_T_15}; // @[Execution.scala 148:64]
  wire [64:0] _data_write_T_16 = _data_write_T_10 | _GEN_11; // @[Execution.scala 148:64]
  wire  _data_write_T_18 = 32'h23 == _mem_wdata_T; // @[Execution.scala 150:39]
  wire [63:0] _data_write_T_20 = _data_write_T_18 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _data_write_T_21 = _data_write_T_20 & data_write_sb; // @[Execution.scala 150:47]
  wire [64:0] _GEN_12 = {{1'd0}, _data_write_T_21}; // @[Execution.scala 149:64]
  wire [64:0] data_write = _data_write_T_16 | _GEN_12; // @[Execution.scala 149:64]
  wire  _data_size_T_4 = _data_write_T_1 | _mem_wdata_T_18; // @[Execution.scala 151:46]
  wire [1:0] _data_size_T_6 = _data_size_T_4 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _data_size_T_15 = _data_write_T_6 | _mem_wdata_T_12 | _mem_wdata_T_36; // @[Execution.scala 152:64]
  wire [1:0] _data_size_T_17 = _data_size_T_15 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _data_size_T_18 = _data_size_T_17 & 2'h2; // @[Execution.scala 152:84]
  wire [1:0] _data_size_T_19 = _data_size_T_6 | _data_size_T_18; // @[Execution.scala 151:94]
  wire  _data_size_T_27 = _data_write_T_12 | _mem_wdata_T_6 | _mem_wdata_T_30; // @[Execution.scala 153:64]
  wire [1:0] _data_size_T_29 = _data_size_T_27 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _data_size_T_30 = _data_size_T_29 & 2'h1; // @[Execution.scala 153:84]
  wire [7:0] _data_strb_T_3 = _data_write_T_1 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _data_strb_T_8 = _data_write_T_6 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _data_strb_T_9 = _data_strb_T_8 & data_strb_sw; // @[Execution.scala 156:47]
  wire [7:0] _data_strb_T_10 = _data_strb_T_3 | _data_strb_T_9; // @[Execution.scala 155:63]
  wire [7:0] _data_strb_T_14 = _data_write_T_12 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _data_strb_T_15 = _data_strb_T_14 & data_strb_sh; // @[Execution.scala 157:47]
  wire [7:0] _data_strb_T_16 = _data_strb_T_10 | _data_strb_T_15; // @[Execution.scala 156:63]
  wire [7:0] _data_strb_T_20 = _data_write_T_18 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _data_strb_T_21 = _data_strb_T_20 & data_strb_sb; // @[Execution.scala 158:47]
  wire [63:0] _ex_wdata_T_1 = io_in_sysop != 4'h0 ? io_csr_rdata : alu_result; // @[Execution.scala 160:48]
  reg [1:0] state; // @[Execution.scala 167:22]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _io_dmem_data_valid_T_1 = state == 2'h0 & data_valid; // @[Execution.scala 188:43]
  assign io_out_valid = io_in_valid; // @[Execution.scala 199:19]
  assign io_out_pc = io_in_pc; // @[Execution.scala 200:19]
  assign io_out_inst = io_in_inst; // @[Execution.scala 201:19]
  assign io_out_wen = io_in_wen; // @[Execution.scala 202:19]
  assign io_out_wdest = io_in_wdest; // @[Execution.scala 203:19]
  assign io_out_wdata = _cmp_ren_T ? mem_wdata : _ex_wdata_T_1; // @[Execution.scala 160:24]
  assign io_out_op1 = io_in_op1; // @[Execution.scala 205:19]
  assign io_out_op2 = io_in_op2; // @[Execution.scala 206:19]
  assign io_out_typew = io_in_typew; // @[Execution.scala 207:19]
  assign io_out_wmem = io_in_wmem; // @[Execution.scala 208:19]
  assign io_out_mem_addr = io_dmem_data_addr; // @[Execution.scala 209:19]
  assign io_out_aluop = io_in_aluop; // @[Execution.scala 211:19]
  assign io_out_loadop = io_in_loadop; // @[Execution.scala 212:19]
  assign io_out_storeop = io_in_storeop; // @[Execution.scala 213:19]
  assign io_out_sysop = io_in_sysop; // @[Execution.scala 214:19]
  assign io_busy = (_io_dmem_data_valid_T_1 | state == 2'h1) & io_in_valid; // @[Execution.scala 195:69]
  assign io_csr_raddr = io_in_inst[31:20]; // @[Execution.scala 75:29]
  assign io_dmem_data_valid = state == 2'h0 & data_valid & io_in_valid; // @[Execution.scala 188:53]
  assign io_dmem_data_req = _cmp_wen_T & _data_valid_T_2; // @[Execution.scala 81:30]
  assign io_dmem_data_addr = alu_result[31:0]; // @[Execution.scala 82:31]
  assign io_dmem_data_size = _data_size_T_19 | _data_size_T_30; // @[Execution.scala 152:94]
  assign io_dmem_data_strb = _data_strb_T_16 | _data_strb_T_21; // @[Execution.scala 157:63]
  assign io_dmem_data_write = data_write[63:0]; // @[Execution.scala 191:23]
  assign io_cmp_ren = io_in_loadop != 7'h0 & (io_dmem_data_addr == 32'h2004000 | io_dmem_data_addr == 32'h200bff8); // @[Execution.scala 64:38]
  assign io_cmp_wen = io_in_storeop != 4'h0 & _cmp_ren_T_3; // @[Execution.scala 65:38]
  assign io_cmp_addr = {{32'd0}, io_dmem_data_addr}; // @[Execution.scala 70:17]
  assign io_cmp_wdata = io_dmem_data_write; // @[Execution.scala 71:17]
  assign io_ex_wdest = io_in_valid ? io_out_wdest : 5'h0; // @[Execution.scala 218:22]
  assign io_ex_result = io_out_wdata; // @[Execution.scala 219:16]
  always @(posedge clock) begin
    if (reset) begin // @[Execution.scala 167:22]
      state <= 2'h0; // @[Execution.scala 167:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (data_valid & io_in_valid) begin // @[Execution.scala 173:33]
        state <= 2'h1; // @[Execution.scala 174:19]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (io_dmem_data_ready) begin // @[Execution.scala 178:27]
        state <= 2'h2; // @[Execution.scala 180:15]
      end
    end else if (_T_3) begin // @[Conditional.scala 39:67]
      state <= 2'h0; // @[Execution.scala 184:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WriteBack(
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_wen,
  input  [4:0]  io_in_wdest,
  input  [63:0] io_in_wdata,
  input  [63:0] io_in_op1,
  input  [31:0] io_in_mem_addr,
  input  [6:0]  io_in_loadop,
  input  [3:0]  io_in_storeop,
  input  [3:0]  io_in_sysop,
  output [31:0] io_pc,
  output [31:0] io_inst,
  output [63:0] io_op1,
  output [3:0]  io_sysop,
  output [6:0]  io_loadop,
  output [3:0]  io_storeop,
  output [31:0] io_mem_addr,
  output        io_wen,
  output [4:0]  io_wdest,
  output [63:0] io_wdata,
  output [4:0]  io_wb_wdest,
  output [63:0] io_wb_result,
  output        io_exc,
  output        io_intr,
  output        io_ready_cmt
);
  wire  _io_intr_T = io_in_sysop == 4'h7; // @[WriteBack.scala 45:23]
  wire  _io_wen_T = ~io_intr; // @[WriteBack.scala 56:30]
  assign io_pc = io_in_pc; // @[WriteBack.scala 48:17]
  assign io_inst = io_in_inst; // @[WriteBack.scala 49:17]
  assign io_op1 = io_in_op1; // @[WriteBack.scala 50:17]
  assign io_sysop = io_in_sysop; // @[WriteBack.scala 51:17]
  assign io_loadop = io_in_loadop; // @[WriteBack.scala 52:17]
  assign io_storeop = io_in_storeop; // @[WriteBack.scala 53:17]
  assign io_mem_addr = io_in_mem_addr; // @[WriteBack.scala 54:17]
  assign io_wen = io_in_wen & ~io_intr & io_in_valid; // @[WriteBack.scala 56:39]
  assign io_wdest = io_in_wdest; // @[WriteBack.scala 57:17]
  assign io_wdata = io_in_wdata; // @[WriteBack.scala 58:17]
  assign io_wb_wdest = io_in_valid ? io_wdest : 5'h0; // @[WriteBack.scala 63:22]
  assign io_wb_result = io_wdata; // @[WriteBack.scala 64:16]
  assign io_exc = io_in_sysop == 4'h4 | io_in_sysop == 4'h5 | _io_intr_T; // @[WriteBack.scala 61:83]
  assign io_intr = io_in_sysop == 4'h7; // @[WriteBack.scala 45:23]
  assign io_ready_cmt = io_in_inst != 32'h0 & _io_wen_T & io_in_valid; // @[WriteBack.scala 59:48]
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_rs1_addr,
  input  [4:0]  io_rs2_addr,
  output [63:0] io_rs1_data,
  output [63:0] io_rs2_data,
  input         io_wen,
  input  [4:0]  io_wdest,
  input  [63:0] io_wdata,
  output [63:0] rf_10
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire  dt_ar_clock; // @[RegFile.scala 25:21]
  wire [7:0] dt_ar_coreid; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_0; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_1; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_2; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_3; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_4; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_5; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_6; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_7; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_8; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_9; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_10; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_11; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_12; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_13; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_14; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_15; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_16; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_17; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_18; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_19; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_20; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_21; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_22; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_23; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_24; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_25; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_26; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_27; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_28; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_29; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_30; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_31; // @[RegFile.scala 25:21]
  reg [63:0] rf__0; // @[RegFile.scala 16:19]
  reg [63:0] rf__1; // @[RegFile.scala 16:19]
  reg [63:0] rf__2; // @[RegFile.scala 16:19]
  reg [63:0] rf__3; // @[RegFile.scala 16:19]
  reg [63:0] rf__4; // @[RegFile.scala 16:19]
  reg [63:0] rf__5; // @[RegFile.scala 16:19]
  reg [63:0] rf__6; // @[RegFile.scala 16:19]
  reg [63:0] rf__7; // @[RegFile.scala 16:19]
  reg [63:0] rf__8; // @[RegFile.scala 16:19]
  reg [63:0] rf__9; // @[RegFile.scala 16:19]
  reg [63:0] rf__10; // @[RegFile.scala 16:19]
  reg [63:0] rf__11; // @[RegFile.scala 16:19]
  reg [63:0] rf__12; // @[RegFile.scala 16:19]
  reg [63:0] rf__13; // @[RegFile.scala 16:19]
  reg [63:0] rf__14; // @[RegFile.scala 16:19]
  reg [63:0] rf__15; // @[RegFile.scala 16:19]
  reg [63:0] rf__16; // @[RegFile.scala 16:19]
  reg [63:0] rf__17; // @[RegFile.scala 16:19]
  reg [63:0] rf__18; // @[RegFile.scala 16:19]
  reg [63:0] rf__19; // @[RegFile.scala 16:19]
  reg [63:0] rf__20; // @[RegFile.scala 16:19]
  reg [63:0] rf__21; // @[RegFile.scala 16:19]
  reg [63:0] rf__22; // @[RegFile.scala 16:19]
  reg [63:0] rf__23; // @[RegFile.scala 16:19]
  reg [63:0] rf__24; // @[RegFile.scala 16:19]
  reg [63:0] rf__25; // @[RegFile.scala 16:19]
  reg [63:0] rf__26; // @[RegFile.scala 16:19]
  reg [63:0] rf__27; // @[RegFile.scala 16:19]
  reg [63:0] rf__28; // @[RegFile.scala 16:19]
  reg [63:0] rf__29; // @[RegFile.scala 16:19]
  reg [63:0] rf__30; // @[RegFile.scala 16:19]
  reg [63:0] rf__31; // @[RegFile.scala 16:19]
  wire [63:0] _GEN_65 = 5'h1 == io_rs1_addr ? rf__1 : rf__0; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_66 = 5'h2 == io_rs1_addr ? rf__2 : _GEN_65; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_67 = 5'h3 == io_rs1_addr ? rf__3 : _GEN_66; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_68 = 5'h4 == io_rs1_addr ? rf__4 : _GEN_67; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_69 = 5'h5 == io_rs1_addr ? rf__5 : _GEN_68; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_70 = 5'h6 == io_rs1_addr ? rf__6 : _GEN_69; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_71 = 5'h7 == io_rs1_addr ? rf__7 : _GEN_70; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_72 = 5'h8 == io_rs1_addr ? rf__8 : _GEN_71; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_73 = 5'h9 == io_rs1_addr ? rf__9 : _GEN_72; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_74 = 5'ha == io_rs1_addr ? rf__10 : _GEN_73; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_75 = 5'hb == io_rs1_addr ? rf__11 : _GEN_74; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_76 = 5'hc == io_rs1_addr ? rf__12 : _GEN_75; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_77 = 5'hd == io_rs1_addr ? rf__13 : _GEN_76; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_78 = 5'he == io_rs1_addr ? rf__14 : _GEN_77; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_79 = 5'hf == io_rs1_addr ? rf__15 : _GEN_78; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_80 = 5'h10 == io_rs1_addr ? rf__16 : _GEN_79; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_81 = 5'h11 == io_rs1_addr ? rf__17 : _GEN_80; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_82 = 5'h12 == io_rs1_addr ? rf__18 : _GEN_81; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_83 = 5'h13 == io_rs1_addr ? rf__19 : _GEN_82; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_84 = 5'h14 == io_rs1_addr ? rf__20 : _GEN_83; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_85 = 5'h15 == io_rs1_addr ? rf__21 : _GEN_84; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_86 = 5'h16 == io_rs1_addr ? rf__22 : _GEN_85; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_87 = 5'h17 == io_rs1_addr ? rf__23 : _GEN_86; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_88 = 5'h18 == io_rs1_addr ? rf__24 : _GEN_87; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_89 = 5'h19 == io_rs1_addr ? rf__25 : _GEN_88; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_90 = 5'h1a == io_rs1_addr ? rf__26 : _GEN_89; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_91 = 5'h1b == io_rs1_addr ? rf__27 : _GEN_90; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_92 = 5'h1c == io_rs1_addr ? rf__28 : _GEN_91; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_93 = 5'h1d == io_rs1_addr ? rf__29 : _GEN_92; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_94 = 5'h1e == io_rs1_addr ? rf__30 : _GEN_93; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_95 = 5'h1f == io_rs1_addr ? rf__31 : _GEN_94; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_97 = 5'h1 == io_rs2_addr ? rf__1 : rf__0; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_98 = 5'h2 == io_rs2_addr ? rf__2 : _GEN_97; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_99 = 5'h3 == io_rs2_addr ? rf__3 : _GEN_98; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_100 = 5'h4 == io_rs2_addr ? rf__4 : _GEN_99; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_101 = 5'h5 == io_rs2_addr ? rf__5 : _GEN_100; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_102 = 5'h6 == io_rs2_addr ? rf__6 : _GEN_101; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_103 = 5'h7 == io_rs2_addr ? rf__7 : _GEN_102; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_104 = 5'h8 == io_rs2_addr ? rf__8 : _GEN_103; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_105 = 5'h9 == io_rs2_addr ? rf__9 : _GEN_104; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_106 = 5'ha == io_rs2_addr ? rf__10 : _GEN_105; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_107 = 5'hb == io_rs2_addr ? rf__11 : _GEN_106; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_108 = 5'hc == io_rs2_addr ? rf__12 : _GEN_107; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_109 = 5'hd == io_rs2_addr ? rf__13 : _GEN_108; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_110 = 5'he == io_rs2_addr ? rf__14 : _GEN_109; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_111 = 5'hf == io_rs2_addr ? rf__15 : _GEN_110; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_112 = 5'h10 == io_rs2_addr ? rf__16 : _GEN_111; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_113 = 5'h11 == io_rs2_addr ? rf__17 : _GEN_112; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_114 = 5'h12 == io_rs2_addr ? rf__18 : _GEN_113; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_115 = 5'h13 == io_rs2_addr ? rf__19 : _GEN_114; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_116 = 5'h14 == io_rs2_addr ? rf__20 : _GEN_115; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_117 = 5'h15 == io_rs2_addr ? rf__21 : _GEN_116; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_118 = 5'h16 == io_rs2_addr ? rf__22 : _GEN_117; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_119 = 5'h17 == io_rs2_addr ? rf__23 : _GEN_118; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_120 = 5'h18 == io_rs2_addr ? rf__24 : _GEN_119; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_121 = 5'h19 == io_rs2_addr ? rf__25 : _GEN_120; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_122 = 5'h1a == io_rs2_addr ? rf__26 : _GEN_121; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_123 = 5'h1b == io_rs2_addr ? rf__27 : _GEN_122; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_124 = 5'h1c == io_rs2_addr ? rf__28 : _GEN_123; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_125 = 5'h1d == io_rs2_addr ? rf__29 : _GEN_124; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_126 = 5'h1e == io_rs2_addr ? rf__30 : _GEN_125; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_127 = 5'h1f == io_rs2_addr ? rf__31 : _GEN_126; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  DifftestArchIntRegState dt_ar ( // @[RegFile.scala 25:21]
    .clock(dt_ar_clock),
    .coreid(dt_ar_coreid),
    .gpr_0(dt_ar_gpr_0),
    .gpr_1(dt_ar_gpr_1),
    .gpr_2(dt_ar_gpr_2),
    .gpr_3(dt_ar_gpr_3),
    .gpr_4(dt_ar_gpr_4),
    .gpr_5(dt_ar_gpr_5),
    .gpr_6(dt_ar_gpr_6),
    .gpr_7(dt_ar_gpr_7),
    .gpr_8(dt_ar_gpr_8),
    .gpr_9(dt_ar_gpr_9),
    .gpr_10(dt_ar_gpr_10),
    .gpr_11(dt_ar_gpr_11),
    .gpr_12(dt_ar_gpr_12),
    .gpr_13(dt_ar_gpr_13),
    .gpr_14(dt_ar_gpr_14),
    .gpr_15(dt_ar_gpr_15),
    .gpr_16(dt_ar_gpr_16),
    .gpr_17(dt_ar_gpr_17),
    .gpr_18(dt_ar_gpr_18),
    .gpr_19(dt_ar_gpr_19),
    .gpr_20(dt_ar_gpr_20),
    .gpr_21(dt_ar_gpr_21),
    .gpr_22(dt_ar_gpr_22),
    .gpr_23(dt_ar_gpr_23),
    .gpr_24(dt_ar_gpr_24),
    .gpr_25(dt_ar_gpr_25),
    .gpr_26(dt_ar_gpr_26),
    .gpr_27(dt_ar_gpr_27),
    .gpr_28(dt_ar_gpr_28),
    .gpr_29(dt_ar_gpr_29),
    .gpr_30(dt_ar_gpr_30),
    .gpr_31(dt_ar_gpr_31)
  );
  assign io_rs1_data = io_rs1_addr != 5'h0 ? _GEN_95 : 64'h0; // @[RegFile.scala 22:21]
  assign io_rs2_data = io_rs2_addr != 5'h0 ? _GEN_127 : 64'h0; // @[RegFile.scala 23:21]
  assign rf_10 = rf__10;
  assign dt_ar_clock = clock; // @[RegFile.scala 26:19]
  assign dt_ar_coreid = 8'h0; // @[RegFile.scala 27:19]
  assign dt_ar_gpr_0 = rf__0; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_1 = rf__1; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_2 = rf__2; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_3 = rf__3; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_4 = rf__4; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_5 = rf__5; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_6 = rf__6; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_7 = rf__7; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_8 = rf__8; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_9 = rf__9; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_10 = rf__10; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_11 = rf__11; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_12 = rf__12; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_13 = rf__13; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_14 = rf__14; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_15 = rf__15; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_16 = rf__16; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_17 = rf__17; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_18 = rf__18; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_19 = rf__19; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_20 = rf__20; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_21 = rf__21; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_22 = rf__22; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_23 = rf__23; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_24 = rf__24; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_25 = rf__25; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_26 = rf__26; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_27 = rf__27; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_28 = rf__28; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_29 = rf__29; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_30 = rf__30; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_31 = rf__31; // @[RegFile.scala 28:19]
  always @(posedge clock) begin
    if (reset) begin // @[RegFile.scala 16:19]
      rf__0 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h0 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__0 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__1 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h1 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__1 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__2 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h2 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__2 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__3 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h3 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__3 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__4 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h4 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__4 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__5 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h5 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__5 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__6 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h6 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__6 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__7 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h7 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__7 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__8 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h8 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__8 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__9 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h9 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__9 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__10 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'ha == io_wdest) begin // @[RegFile.scala 19:18]
        rf__10 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__11 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'hb == io_wdest) begin // @[RegFile.scala 19:18]
        rf__11 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__12 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'hc == io_wdest) begin // @[RegFile.scala 19:18]
        rf__12 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__13 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'hd == io_wdest) begin // @[RegFile.scala 19:18]
        rf__13 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__14 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'he == io_wdest) begin // @[RegFile.scala 19:18]
        rf__14 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__15 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'hf == io_wdest) begin // @[RegFile.scala 19:18]
        rf__15 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__16 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h10 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__16 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__17 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h11 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__17 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__18 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h12 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__18 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__19 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h13 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__19 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__20 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h14 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__20 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__21 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h15 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__21 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__22 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h16 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__22 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__23 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h17 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__23 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__24 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h18 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__24 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__25 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h19 == io_wdest) begin // @[RegFile.scala 19:18]
        rf__25 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__26 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h1a == io_wdest) begin // @[RegFile.scala 19:18]
        rf__26 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__27 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h1b == io_wdest) begin // @[RegFile.scala 19:18]
        rf__27 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__28 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h1c == io_wdest) begin // @[RegFile.scala 19:18]
        rf__28 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__29 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h1d == io_wdest) begin // @[RegFile.scala 19:18]
        rf__29 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__30 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h1e == io_wdest) begin // @[RegFile.scala 19:18]
        rf__30 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__31 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_wen & io_wdest != 5'h0) begin // @[RegFile.scala 18:39]
      if (5'h1f == io_wdest) begin // @[RegFile.scala 19:18]
        rf__31 <= io_wdata; // @[RegFile.scala 19:18]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rf__0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  rf__1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf__2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf__3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf__4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf__5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf__6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf__7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf__8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf__9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf__10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf__11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf__12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf__13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf__14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf__15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf__16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf__17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf__18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf__19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf__20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf__21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf__22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf__23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf__24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf__25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf__26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf__27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf__28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf__29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf__30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  rf__31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Csr(
  input         clock,
  input         reset,
  input  [63:0] io_in1,
  input  [31:0] io_pc,
  input  [31:0] io_inst,
  input  [11:0] io_raddr,
  input  [3:0]  io_sysop,
  input         io_exc,
  output [63:0] io_csr_rdata,
  output [63:0] io_mstatus,
  output [63:0] io_mie,
  output [63:0] io_mtvec,
  output [63:0] io_mepc
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  dt_cs_clock; // @[Csr.scala 133:21]
  wire [7:0] dt_cs_coreid; // @[Csr.scala 133:21]
  wire [1:0] dt_cs_priviledgeMode; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_mstatus; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_sstatus; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_mepc; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_sepc; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_mtval; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_stval; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_mtvec; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_stvec; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_mcause; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_scause; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_satp; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_mip; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_mie; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_mscratch; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_sscratch; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_mideleg; // @[Csr.scala 133:21]
  wire [63:0] dt_cs_medeleg; // @[Csr.scala 133:21]
  wire [4:0] in2_lo = io_inst[19:15]; // @[Csr.scala 25:39]
  wire [63:0] in2 = {59'h0,in2_lo}; // @[Cat.scala 30:58]
  wire  _csr_rw_T = io_sysop == 4'h1; // @[Csr.scala 27:23]
  wire  _csr_rw_T_1 = io_sysop == 4'h2; // @[Csr.scala 28:23]
  wire  _csr_rw_T_2 = io_sysop == 4'h1 | _csr_rw_T_1; // @[Csr.scala 27:46]
  wire  _csr_rw_T_4 = _csr_rw_T_2 | _csr_rw_T; // @[Csr.scala 28:46]
  wire  _csr_rw_T_5 = io_sysop == 4'h8; // @[Csr.scala 30:23]
  wire  _csr_rw_T_6 = _csr_rw_T_4 | _csr_rw_T_5; // @[Csr.scala 29:46]
  wire  _csr_rw_T_7 = io_sysop == 4'h9; // @[Csr.scala 31:23]
  wire  csr_rw = _csr_rw_T_6 | _csr_rw_T_7; // @[Csr.scala 30:46]
  reg [63:0] mstatus; // @[Csr.scala 34:26]
  reg [63:0] mie; // @[Csr.scala 35:26]
  reg [63:0] mtvec; // @[Csr.scala 37:26]
  reg [63:0] mscratch; // @[Csr.scala 38:26]
  reg [63:0] mepc; // @[Csr.scala 39:26]
  reg [63:0] mcause; // @[Csr.scala 40:26]
  reg [63:0] mcycle; // @[Csr.scala 41:26]
  wire [50:0] mstatus_hi_hi_hi = mstatus[63:13]; // @[Csr.scala 48:27]
  wire [2:0] mstatus_hi_lo_hi = mstatus[10:8]; // @[Csr.scala 48:57]
  wire  mstatus_hi_lo_lo = mstatus[3]; // @[Csr.scala 48:72]
  wire [2:0] mstatus_lo_hi_hi = mstatus[6:4]; // @[Csr.scala 48:84]
  wire [2:0] mstatus_lo_lo = mstatus[2:0]; // @[Csr.scala 48:104]
  wire [63:0] _mstatus_T = {mstatus_hi_hi_hi,2'h3,mstatus_hi_lo_hi,mstatus_hi_lo_lo,mstatus_lo_hi_hi,1'h0,mstatus_lo_lo}
    ; // @[Cat.scala 30:58]
  wire [63:0] _GEN_0 = io_sysop == 4'h4 & io_exc ? {{32'd0}, io_pc} : mepc; // @[Csr.scala 45:47 Csr.scala 46:10 Csr.scala 39:26]
  wire [63:0] _GEN_1 = io_sysop == 4'h4 & io_exc ? 64'hb : mcause; // @[Csr.scala 45:47 Csr.scala 47:12 Csr.scala 40:26]
  wire [63:0] _GEN_2 = io_sysop == 4'h4 & io_exc ? _mstatus_T : mstatus; // @[Csr.scala 45:47 Csr.scala 48:13 Csr.scala 34:26]
  wire  mstatus_lo_hi_lo = mstatus[7]; // @[Csr.scala 53:92]
  wire [63:0] _mstatus_T_1 = {mstatus_hi_hi_hi,2'h0,mstatus_hi_lo_hi,1'h1,mstatus_lo_hi_hi,mstatus_lo_hi_lo,
    mstatus_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_3 = io_sysop == 4'h5 & io_exc ? _mstatus_T_1 : _GEN_2; // @[Csr.scala 52:46 Csr.scala 53:13]
  wire [63:0] _GEN_4 = io_sysop == 4'h7 & io_exc ? {{32'd0}, io_pc} : _GEN_0; // @[Csr.scala 57:45 Csr.scala 58:10]
  wire [63:0] _GEN_5 = io_sysop == 4'h7 & io_exc ? 64'h8000000000000007 : _GEN_1; // @[Csr.scala 57:45 Csr.scala 59:12]
  wire [63:0] _GEN_6 = io_sysop == 4'h7 & io_exc ? _mstatus_T : _GEN_3; // @[Csr.scala 57:45 Csr.scala 60:13]
  wire [11:0] waddr = io_inst[31:20]; // @[Csr.scala 64:22]
  wire [63:0] _op1_T_1 = 12'h300 == waddr ? mstatus : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _op1_T_3 = 12'h342 == waddr ? mcause : _op1_T_1; // @[Mux.scala 80:57]
  wire [63:0] _op1_T_5 = 12'h304 == waddr ? mie : _op1_T_3; // @[Mux.scala 80:57]
  wire [63:0] _op1_T_7 = 12'h305 == waddr ? mtvec : _op1_T_5; // @[Mux.scala 80:57]
  wire [63:0] _op1_T_9 = 12'h340 == waddr ? mscratch : _op1_T_7; // @[Mux.scala 80:57]
  wire [63:0] _op1_T_11 = 12'h341 == waddr ? mepc : _op1_T_9; // @[Mux.scala 80:57]
  wire [63:0] _op1_T_13 = 12'h344 == waddr ? 64'h0 : _op1_T_11; // @[Mux.scala 80:57]
  wire [63:0] _op1_T_15 = 12'hb00 == waddr ? mcycle : _op1_T_13; // @[Mux.scala 80:57]
  wire [63:0] op1 = 12'hb02 == waddr ? 64'h0 : _op1_T_15; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_1 = 12'h300 == io_raddr ? mstatus : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_3 = 12'h342 == io_raddr ? mcause : _rdata_T_1; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_5 = 12'h304 == io_raddr ? mie : _rdata_T_3; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_7 = 12'h305 == io_raddr ? mtvec : _rdata_T_5; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_9 = 12'h340 == io_raddr ? mscratch : _rdata_T_7; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_11 = 12'h341 == io_raddr ? mepc : _rdata_T_9; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_13 = 12'h344 == io_raddr ? 64'h0 : _rdata_T_11; // @[Mux.scala 80:57]
  wire [63:0] _rdata_T_15 = 12'hb00 == io_raddr ? mcycle : _rdata_T_13; // @[Mux.scala 80:57]
  wire [63:0] _wdata_T = op1 | io_in1; // @[Csr.scala 93:43]
  wire [63:0] _wdata_T_1 = ~io_in1; // @[Csr.scala 94:45]
  wire [63:0] _wdata_T_2 = op1 & _wdata_T_1; // @[Csr.scala 94:43]
  wire [63:0] _wdata_T_3 = op1 | in2; // @[Csr.scala 95:43]
  wire [63:0] _wdata_T_4 = ~in2; // @[Csr.scala 96:45]
  wire [63:0] _wdata_T_5 = op1 & _wdata_T_4; // @[Csr.scala 96:43]
  wire [63:0] _wdata_T_7 = 4'h1 == io_sysop ? io_in1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _wdata_T_9 = 4'h2 == io_sysop ? _wdata_T : _wdata_T_7; // @[Mux.scala 80:57]
  wire [63:0] _wdata_T_11 = 4'h3 == io_sysop ? _wdata_T_2 : _wdata_T_9; // @[Mux.scala 80:57]
  wire [63:0] _wdata_T_13 = 4'h8 == io_sysop ? _wdata_T_3 : _wdata_T_11; // @[Mux.scala 80:57]
  wire [63:0] wdata = 4'h9 == io_sysop ? _wdata_T_5 : _wdata_T_13; // @[Mux.scala 80:57]
  wire [63:0] _mcycle_T_1 = mcycle + 64'h1; // @[Csr.scala 100:20]
  wire  mstatus_hi_3 = wdata[16] & wdata[15] | wdata[14] & wdata[13]; // @[Csr.scala 116:46]
  wire [62:0] mstatus_lo_3 = wdata[62:0]; // @[Csr.scala 116:79]
  wire [63:0] _mstatus_T_9 = {mstatus_hi_3,mstatus_lo_3}; // @[Cat.scala 30:58]
  DifftestCSRState dt_cs ( // @[Csr.scala 133:21]
    .clock(dt_cs_clock),
    .coreid(dt_cs_coreid),
    .priviledgeMode(dt_cs_priviledgeMode),
    .mstatus(dt_cs_mstatus),
    .sstatus(dt_cs_sstatus),
    .mepc(dt_cs_mepc),
    .sepc(dt_cs_sepc),
    .mtval(dt_cs_mtval),
    .stval(dt_cs_stval),
    .mtvec(dt_cs_mtvec),
    .stvec(dt_cs_stvec),
    .mcause(dt_cs_mcause),
    .scause(dt_cs_scause),
    .satp(dt_cs_satp),
    .mip(dt_cs_mip),
    .mie(dt_cs_mie),
    .mscratch(dt_cs_mscratch),
    .sscratch(dt_cs_sscratch),
    .mideleg(dt_cs_mideleg),
    .medeleg(dt_cs_medeleg)
  );
  assign io_csr_rdata = 12'hb02 == io_raddr ? 64'h0 : _rdata_T_15; // @[Mux.scala 80:57]
  assign io_mstatus = mstatus; // @[Csr.scala 127:17]
  assign io_mie = mie; // @[Csr.scala 128:17]
  assign io_mtvec = mtvec; // @[Csr.scala 129:17]
  assign io_mepc = mepc; // @[Csr.scala 130:17]
  assign dt_cs_clock = clock; // @[Csr.scala 134:27]
  assign dt_cs_coreid = 8'h0; // @[Csr.scala 135:27]
  assign dt_cs_priviledgeMode = 2'h3; // @[Csr.scala 136:27]
  assign dt_cs_mstatus = mstatus; // @[Csr.scala 137:27]
  assign dt_cs_sstatus = mstatus & 64'h80000003000de122; // @[Csr.scala 138:38]
  assign dt_cs_mepc = mepc; // @[Csr.scala 139:27]
  assign dt_cs_sepc = 64'h0; // @[Csr.scala 140:27]
  assign dt_cs_mtval = 64'h0; // @[Csr.scala 141:27]
  assign dt_cs_stval = 64'h0; // @[Csr.scala 142:27]
  assign dt_cs_mtvec = mtvec; // @[Csr.scala 143:27]
  assign dt_cs_stvec = 64'h0; // @[Csr.scala 144:27]
  assign dt_cs_mcause = mcause; // @[Csr.scala 145:27]
  assign dt_cs_scause = 64'h0; // @[Csr.scala 146:27]
  assign dt_cs_satp = 64'h0; // @[Csr.scala 147:27]
  assign dt_cs_mip = 64'h0; // @[Csr.scala 148:27]
  assign dt_cs_mie = mie; // @[Csr.scala 149:27]
  assign dt_cs_mscratch = mscratch; // @[Csr.scala 150:27]
  assign dt_cs_sscratch = 64'h0; // @[Csr.scala 151:27]
  assign dt_cs_mideleg = 64'h0; // @[Csr.scala 152:27]
  assign dt_cs_medeleg = 64'h0; // @[Csr.scala 153:27]
  always @(posedge clock) begin
    if (reset) begin // @[Csr.scala 34:26]
      mstatus <= 64'h1800; // @[Csr.scala 34:26]
    end else if (csr_rw) begin // @[Csr.scala 102:13]
      if (waddr == 12'h300) begin // @[Csr.scala 115:34]
        mstatus <= _mstatus_T_9; // @[Csr.scala 116:15]
      end else begin
        mstatus <= _GEN_6;
      end
    end else begin
      mstatus <= _GEN_6;
    end
    if (reset) begin // @[Csr.scala 35:26]
      mie <= 64'h0; // @[Csr.scala 35:26]
    end else if (csr_rw) begin // @[Csr.scala 102:13]
      if (waddr == 12'h304) begin // @[Csr.scala 118:30]
        if (4'h9 == io_sysop) begin // @[Mux.scala 80:57]
          mie <= _wdata_T_5;
        end else begin
          mie <= _wdata_T_13;
        end
      end
    end
    if (reset) begin // @[Csr.scala 37:26]
      mtvec <= 64'h0; // @[Csr.scala 37:26]
    end else if (csr_rw) begin // @[Csr.scala 102:13]
      if (waddr == 12'h305) begin // @[Csr.scala 106:32]
        if (4'h9 == io_sysop) begin // @[Mux.scala 80:57]
          mtvec <= _wdata_T_5;
        end else begin
          mtvec <= _wdata_T_13;
        end
      end
    end
    if (reset) begin // @[Csr.scala 38:26]
      mscratch <= 64'h0; // @[Csr.scala 38:26]
    end else if (csr_rw) begin // @[Csr.scala 102:13]
      if (waddr == 12'h340) begin // @[Csr.scala 121:35]
        if (4'h9 == io_sysop) begin // @[Mux.scala 80:57]
          mscratch <= _wdata_T_5;
        end else begin
          mscratch <= _wdata_T_13;
        end
      end
    end
    if (reset) begin // @[Csr.scala 39:26]
      mepc <= 64'h0; // @[Csr.scala 39:26]
    end else if (csr_rw) begin // @[Csr.scala 102:13]
      if (waddr == 12'h341) begin // @[Csr.scala 109:31]
        if (4'h9 == io_sysop) begin // @[Mux.scala 80:57]
          mepc <= _wdata_T_5;
        end else begin
          mepc <= _wdata_T_13;
        end
      end else begin
        mepc <= _GEN_4;
      end
    end else begin
      mepc <= _GEN_4;
    end
    if (reset) begin // @[Csr.scala 40:26]
      mcause <= 64'h0; // @[Csr.scala 40:26]
    end else if (csr_rw) begin // @[Csr.scala 102:13]
      if (waddr == 12'h342) begin // @[Csr.scala 112:33]
        if (4'h9 == io_sysop) begin // @[Mux.scala 80:57]
          mcause <= _wdata_T_5;
        end else begin
          mcause <= _wdata_T_13;
        end
      end else begin
        mcause <= _GEN_5;
      end
    end else begin
      mcause <= _GEN_5;
    end
    if (reset) begin // @[Csr.scala 41:26]
      mcycle <= 64'h0; // @[Csr.scala 41:26]
    end else if (csr_rw) begin // @[Csr.scala 102:13]
      if (waddr == 12'hb00) begin // @[Csr.scala 103:33]
        if (4'h9 == io_sysop) begin // @[Mux.scala 80:57]
          mcycle <= _wdata_T_5;
        end else begin
          mcycle <= _wdata_T_13;
        end
      end else begin
        mcycle <= _mcycle_T_1; // @[Csr.scala 100:10]
      end
    end else begin
      mcycle <= _mcycle_T_1; // @[Csr.scala 100:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mstatus = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mie = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mtvec = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mscratch = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mepc = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mcause = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mcycle = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Clint(
  input         clock,
  input         reset,
  input  [63:0] io_mstatus,
  input  [63:0] io_mie,
  input         io_exc,
  input         io_cmp_ren,
  input         io_cmp_wen,
  input  [63:0] io_cmp_addr,
  input  [63:0] io_cmp_wdata,
  output [63:0] io_cmp_rdata,
  output        io_time_int
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[Clint.scala 28:26]
  reg [63:0] mtimecmp; // @[Clint.scala 29:26]
  wire [63:0] _mtime_T_1 = mtime + 64'h1; // @[Clint.scala 31:18]
  wire [63:0] _io_cmp_rdata_T_1 = io_cmp_addr == 64'h200bff8 ? mtime : mtimecmp; // @[Clint.scala 38:35]
  assign io_cmp_rdata = io_cmp_ren ? _io_cmp_rdata_T_1 : 64'h0; // @[Clint.scala 38:22]
  assign io_time_int = mtime >= mtimecmp & io_mstatus[3] & io_mie[7] & ~io_exc; // @[Clint.scala 36:77]
  always @(posedge clock) begin
    if (reset) begin // @[Clint.scala 28:26]
      mtime <= 64'h0; // @[Clint.scala 28:26]
    end else begin
      mtime <= _mtime_T_1; // @[Clint.scala 31:9]
    end
    if (reset) begin // @[Clint.scala 29:26]
      mtimecmp <= 64'h0; // @[Clint.scala 29:26]
    end else if (io_cmp_wen) begin // @[Clint.scala 32:18]
      mtimecmp <= io_cmp_wdata; // @[Clint.scala 33:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core(
  input         clock,
  input         reset,
  output        io_imem_inst_valid,
  input         io_imem_inst_ready,
  output [31:0] io_imem_inst_addr,
  input  [31:0] io_imem_inst_read,
  output        io_dmem_data_valid,
  input         io_dmem_data_ready,
  output        io_dmem_data_req,
  output [31:0] io_dmem_data_addr,
  output [1:0]  io_dmem_data_size,
  output [7:0]  io_dmem_data_strb,
  input  [63:0] io_dmem_data_read,
  output [63:0] io_dmem_data_write
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  fetch_clock; // @[Core.scala 13:21]
  wire  fetch_reset; // @[Core.scala 13:21]
  wire  fetch_io_imem_inst_valid; // @[Core.scala 13:21]
  wire  fetch_io_imem_inst_ready; // @[Core.scala 13:21]
  wire [31:0] fetch_io_imem_inst_addr; // @[Core.scala 13:21]
  wire [31:0] fetch_io_imem_inst_read; // @[Core.scala 13:21]
  wire  fetch_io_jmp_packet_valid; // @[Core.scala 13:21]
  wire [31:0] fetch_io_jmp_packet_inst_pc; // @[Core.scala 13:21]
  wire  fetch_io_jmp_packet_jmp; // @[Core.scala 13:21]
  wire [31:0] fetch_io_jmp_packet_jmp_pc; // @[Core.scala 13:21]
  wire  fetch_io_jmp_packet_mis; // @[Core.scala 13:21]
  wire  fetch_io_stall; // @[Core.scala 13:21]
  wire  fetch_io_out_valid; // @[Core.scala 13:21]
  wire [31:0] fetch_io_out_pc; // @[Core.scala 13:21]
  wire [31:0] fetch_io_out_inst; // @[Core.scala 13:21]
  wire  fetch_io_out_bp_taken; // @[Core.scala 13:21]
  wire [31:0] fetch_io_out_bp_targer; // @[Core.scala 13:21]
  wire  reg_if_id_clock; // @[Core.scala 14:25]
  wire  reg_if_id_reset; // @[Core.scala 14:25]
  wire  reg_if_id_io_in_valid; // @[Core.scala 14:25]
  wire [31:0] reg_if_id_io_in_pc; // @[Core.scala 14:25]
  wire [31:0] reg_if_id_io_in_inst; // @[Core.scala 14:25]
  wire  reg_if_id_io_in_wen; // @[Core.scala 14:25]
  wire [4:0] reg_if_id_io_in_wdest; // @[Core.scala 14:25]
  wire [63:0] reg_if_id_io_in_wdata; // @[Core.scala 14:25]
  wire [63:0] reg_if_id_io_in_op1; // @[Core.scala 14:25]
  wire [63:0] reg_if_id_io_in_op2; // @[Core.scala 14:25]
  wire  reg_if_id_io_in_typew; // @[Core.scala 14:25]
  wire [63:0] reg_if_id_io_in_wmem; // @[Core.scala 14:25]
  wire [31:0] reg_if_id_io_in_mem_addr; // @[Core.scala 14:25]
  wire [11:0] reg_if_id_io_in_aluop; // @[Core.scala 14:25]
  wire [6:0] reg_if_id_io_in_loadop; // @[Core.scala 14:25]
  wire [3:0] reg_if_id_io_in_storeop; // @[Core.scala 14:25]
  wire [3:0] reg_if_id_io_in_sysop; // @[Core.scala 14:25]
  wire  reg_if_id_io_in_bp_taken; // @[Core.scala 14:25]
  wire [31:0] reg_if_id_io_in_bp_targer; // @[Core.scala 14:25]
  wire  reg_if_id_io_out_valid; // @[Core.scala 14:25]
  wire [31:0] reg_if_id_io_out_pc; // @[Core.scala 14:25]
  wire [31:0] reg_if_id_io_out_inst; // @[Core.scala 14:25]
  wire  reg_if_id_io_out_wen; // @[Core.scala 14:25]
  wire [4:0] reg_if_id_io_out_wdest; // @[Core.scala 14:25]
  wire [63:0] reg_if_id_io_out_wdata; // @[Core.scala 14:25]
  wire [63:0] reg_if_id_io_out_op1; // @[Core.scala 14:25]
  wire [63:0] reg_if_id_io_out_op2; // @[Core.scala 14:25]
  wire  reg_if_id_io_out_typew; // @[Core.scala 14:25]
  wire [63:0] reg_if_id_io_out_wmem; // @[Core.scala 14:25]
  wire [31:0] reg_if_id_io_out_mem_addr; // @[Core.scala 14:25]
  wire [11:0] reg_if_id_io_out_aluop; // @[Core.scala 14:25]
  wire [6:0] reg_if_id_io_out_loadop; // @[Core.scala 14:25]
  wire [3:0] reg_if_id_io_out_storeop; // @[Core.scala 14:25]
  wire [3:0] reg_if_id_io_out_sysop; // @[Core.scala 14:25]
  wire  reg_if_id_io_out_bp_taken; // @[Core.scala 14:25]
  wire [31:0] reg_if_id_io_out_bp_targer; // @[Core.scala 14:25]
  wire  reg_if_id_io_stall; // @[Core.scala 14:25]
  wire [4:0] decode_io_rs1_addr; // @[Core.scala 15:22]
  wire [4:0] decode_io_rs2_addr; // @[Core.scala 15:22]
  wire [63:0] decode_io_rs1_data; // @[Core.scala 15:22]
  wire [63:0] decode_io_rs2_data; // @[Core.scala 15:22]
  wire  decode_io_in_valid; // @[Core.scala 15:22]
  wire [31:0] decode_io_in_pc; // @[Core.scala 15:22]
  wire [31:0] decode_io_in_inst; // @[Core.scala 15:22]
  wire  decode_io_in_bp_taken; // @[Core.scala 15:22]
  wire [31:0] decode_io_in_bp_targer; // @[Core.scala 15:22]
  wire  decode_io_out_valid; // @[Core.scala 15:22]
  wire [31:0] decode_io_out_pc; // @[Core.scala 15:22]
  wire [31:0] decode_io_out_inst; // @[Core.scala 15:22]
  wire  decode_io_out_wen; // @[Core.scala 15:22]
  wire [4:0] decode_io_out_wdest; // @[Core.scala 15:22]
  wire [63:0] decode_io_out_op1; // @[Core.scala 15:22]
  wire [63:0] decode_io_out_op2; // @[Core.scala 15:22]
  wire  decode_io_out_typew; // @[Core.scala 15:22]
  wire [63:0] decode_io_out_wmem; // @[Core.scala 15:22]
  wire [11:0] decode_io_out_aluop; // @[Core.scala 15:22]
  wire [6:0] decode_io_out_loadop; // @[Core.scala 15:22]
  wire [3:0] decode_io_out_storeop; // @[Core.scala 15:22]
  wire [3:0] decode_io_out_sysop; // @[Core.scala 15:22]
  wire  decode_io_jmp_packet_valid; // @[Core.scala 15:22]
  wire [31:0] decode_io_jmp_packet_inst_pc; // @[Core.scala 15:22]
  wire  decode_io_jmp_packet_jmp; // @[Core.scala 15:22]
  wire [31:0] decode_io_jmp_packet_jmp_pc; // @[Core.scala 15:22]
  wire  decode_io_jmp_packet_mis; // @[Core.scala 15:22]
  wire  decode_io_stall; // @[Core.scala 15:22]
  wire [63:0] decode_io_mtvec; // @[Core.scala 15:22]
  wire [63:0] decode_io_mepc; // @[Core.scala 15:22]
  wire  decode_io_time_int; // @[Core.scala 15:22]
  wire [4:0] decode_io_ex_wdest; // @[Core.scala 15:22]
  wire [4:0] decode_io_wb_wdest; // @[Core.scala 15:22]
  wire [63:0] decode_io_ex_result; // @[Core.scala 15:22]
  wire [63:0] decode_io_wb_result; // @[Core.scala 15:22]
  wire  reg_id_ex_clock; // @[Core.scala 16:25]
  wire  reg_id_ex_reset; // @[Core.scala 16:25]
  wire  reg_id_ex_io_in_valid; // @[Core.scala 16:25]
  wire [31:0] reg_id_ex_io_in_pc; // @[Core.scala 16:25]
  wire [31:0] reg_id_ex_io_in_inst; // @[Core.scala 16:25]
  wire  reg_id_ex_io_in_wen; // @[Core.scala 16:25]
  wire [4:0] reg_id_ex_io_in_wdest; // @[Core.scala 16:25]
  wire [63:0] reg_id_ex_io_in_wdata; // @[Core.scala 16:25]
  wire [63:0] reg_id_ex_io_in_op1; // @[Core.scala 16:25]
  wire [63:0] reg_id_ex_io_in_op2; // @[Core.scala 16:25]
  wire  reg_id_ex_io_in_typew; // @[Core.scala 16:25]
  wire [63:0] reg_id_ex_io_in_wmem; // @[Core.scala 16:25]
  wire [31:0] reg_id_ex_io_in_mem_addr; // @[Core.scala 16:25]
  wire [11:0] reg_id_ex_io_in_aluop; // @[Core.scala 16:25]
  wire [6:0] reg_id_ex_io_in_loadop; // @[Core.scala 16:25]
  wire [3:0] reg_id_ex_io_in_storeop; // @[Core.scala 16:25]
  wire [3:0] reg_id_ex_io_in_sysop; // @[Core.scala 16:25]
  wire  reg_id_ex_io_in_bp_taken; // @[Core.scala 16:25]
  wire [31:0] reg_id_ex_io_in_bp_targer; // @[Core.scala 16:25]
  wire  reg_id_ex_io_out_valid; // @[Core.scala 16:25]
  wire [31:0] reg_id_ex_io_out_pc; // @[Core.scala 16:25]
  wire [31:0] reg_id_ex_io_out_inst; // @[Core.scala 16:25]
  wire  reg_id_ex_io_out_wen; // @[Core.scala 16:25]
  wire [4:0] reg_id_ex_io_out_wdest; // @[Core.scala 16:25]
  wire [63:0] reg_id_ex_io_out_wdata; // @[Core.scala 16:25]
  wire [63:0] reg_id_ex_io_out_op1; // @[Core.scala 16:25]
  wire [63:0] reg_id_ex_io_out_op2; // @[Core.scala 16:25]
  wire  reg_id_ex_io_out_typew; // @[Core.scala 16:25]
  wire [63:0] reg_id_ex_io_out_wmem; // @[Core.scala 16:25]
  wire [31:0] reg_id_ex_io_out_mem_addr; // @[Core.scala 16:25]
  wire [11:0] reg_id_ex_io_out_aluop; // @[Core.scala 16:25]
  wire [6:0] reg_id_ex_io_out_loadop; // @[Core.scala 16:25]
  wire [3:0] reg_id_ex_io_out_storeop; // @[Core.scala 16:25]
  wire [3:0] reg_id_ex_io_out_sysop; // @[Core.scala 16:25]
  wire  reg_id_ex_io_out_bp_taken; // @[Core.scala 16:25]
  wire [31:0] reg_id_ex_io_out_bp_targer; // @[Core.scala 16:25]
  wire  reg_id_ex_io_stall; // @[Core.scala 16:25]
  wire  execution_clock; // @[Core.scala 17:25]
  wire  execution_reset; // @[Core.scala 17:25]
  wire  execution_io_in_valid; // @[Core.scala 17:25]
  wire [31:0] execution_io_in_pc; // @[Core.scala 17:25]
  wire [31:0] execution_io_in_inst; // @[Core.scala 17:25]
  wire  execution_io_in_wen; // @[Core.scala 17:25]
  wire [4:0] execution_io_in_wdest; // @[Core.scala 17:25]
  wire [63:0] execution_io_in_op1; // @[Core.scala 17:25]
  wire [63:0] execution_io_in_op2; // @[Core.scala 17:25]
  wire  execution_io_in_typew; // @[Core.scala 17:25]
  wire [63:0] execution_io_in_wmem; // @[Core.scala 17:25]
  wire [11:0] execution_io_in_aluop; // @[Core.scala 17:25]
  wire [6:0] execution_io_in_loadop; // @[Core.scala 17:25]
  wire [3:0] execution_io_in_storeop; // @[Core.scala 17:25]
  wire [3:0] execution_io_in_sysop; // @[Core.scala 17:25]
  wire  execution_io_out_valid; // @[Core.scala 17:25]
  wire [31:0] execution_io_out_pc; // @[Core.scala 17:25]
  wire [31:0] execution_io_out_inst; // @[Core.scala 17:25]
  wire  execution_io_out_wen; // @[Core.scala 17:25]
  wire [4:0] execution_io_out_wdest; // @[Core.scala 17:25]
  wire [63:0] execution_io_out_wdata; // @[Core.scala 17:25]
  wire [63:0] execution_io_out_op1; // @[Core.scala 17:25]
  wire [63:0] execution_io_out_op2; // @[Core.scala 17:25]
  wire  execution_io_out_typew; // @[Core.scala 17:25]
  wire [63:0] execution_io_out_wmem; // @[Core.scala 17:25]
  wire [31:0] execution_io_out_mem_addr; // @[Core.scala 17:25]
  wire [11:0] execution_io_out_aluop; // @[Core.scala 17:25]
  wire [6:0] execution_io_out_loadop; // @[Core.scala 17:25]
  wire [3:0] execution_io_out_storeop; // @[Core.scala 17:25]
  wire [3:0] execution_io_out_sysop; // @[Core.scala 17:25]
  wire  execution_io_busy; // @[Core.scala 17:25]
  wire [11:0] execution_io_csr_raddr; // @[Core.scala 17:25]
  wire [63:0] execution_io_csr_rdata; // @[Core.scala 17:25]
  wire  execution_io_dmem_data_valid; // @[Core.scala 17:25]
  wire  execution_io_dmem_data_ready; // @[Core.scala 17:25]
  wire  execution_io_dmem_data_req; // @[Core.scala 17:25]
  wire [31:0] execution_io_dmem_data_addr; // @[Core.scala 17:25]
  wire [1:0] execution_io_dmem_data_size; // @[Core.scala 17:25]
  wire [7:0] execution_io_dmem_data_strb; // @[Core.scala 17:25]
  wire [63:0] execution_io_dmem_data_read; // @[Core.scala 17:25]
  wire [63:0] execution_io_dmem_data_write; // @[Core.scala 17:25]
  wire  execution_io_cmp_ren; // @[Core.scala 17:25]
  wire  execution_io_cmp_wen; // @[Core.scala 17:25]
  wire [63:0] execution_io_cmp_addr; // @[Core.scala 17:25]
  wire [63:0] execution_io_cmp_wdata; // @[Core.scala 17:25]
  wire [63:0] execution_io_cmp_rdata; // @[Core.scala 17:25]
  wire [4:0] execution_io_ex_wdest; // @[Core.scala 17:25]
  wire [63:0] execution_io_ex_result; // @[Core.scala 17:25]
  wire  reg_ex_wb_clock; // @[Core.scala 18:25]
  wire  reg_ex_wb_reset; // @[Core.scala 18:25]
  wire  reg_ex_wb_io_in_valid; // @[Core.scala 18:25]
  wire [31:0] reg_ex_wb_io_in_pc; // @[Core.scala 18:25]
  wire [31:0] reg_ex_wb_io_in_inst; // @[Core.scala 18:25]
  wire  reg_ex_wb_io_in_wen; // @[Core.scala 18:25]
  wire [4:0] reg_ex_wb_io_in_wdest; // @[Core.scala 18:25]
  wire [63:0] reg_ex_wb_io_in_wdata; // @[Core.scala 18:25]
  wire [63:0] reg_ex_wb_io_in_op1; // @[Core.scala 18:25]
  wire [63:0] reg_ex_wb_io_in_op2; // @[Core.scala 18:25]
  wire  reg_ex_wb_io_in_typew; // @[Core.scala 18:25]
  wire [63:0] reg_ex_wb_io_in_wmem; // @[Core.scala 18:25]
  wire [31:0] reg_ex_wb_io_in_mem_addr; // @[Core.scala 18:25]
  wire [11:0] reg_ex_wb_io_in_aluop; // @[Core.scala 18:25]
  wire [6:0] reg_ex_wb_io_in_loadop; // @[Core.scala 18:25]
  wire [3:0] reg_ex_wb_io_in_storeop; // @[Core.scala 18:25]
  wire [3:0] reg_ex_wb_io_in_sysop; // @[Core.scala 18:25]
  wire  reg_ex_wb_io_in_bp_taken; // @[Core.scala 18:25]
  wire [31:0] reg_ex_wb_io_in_bp_targer; // @[Core.scala 18:25]
  wire  reg_ex_wb_io_out_valid; // @[Core.scala 18:25]
  wire [31:0] reg_ex_wb_io_out_pc; // @[Core.scala 18:25]
  wire [31:0] reg_ex_wb_io_out_inst; // @[Core.scala 18:25]
  wire  reg_ex_wb_io_out_wen; // @[Core.scala 18:25]
  wire [4:0] reg_ex_wb_io_out_wdest; // @[Core.scala 18:25]
  wire [63:0] reg_ex_wb_io_out_wdata; // @[Core.scala 18:25]
  wire [63:0] reg_ex_wb_io_out_op1; // @[Core.scala 18:25]
  wire [63:0] reg_ex_wb_io_out_op2; // @[Core.scala 18:25]
  wire  reg_ex_wb_io_out_typew; // @[Core.scala 18:25]
  wire [63:0] reg_ex_wb_io_out_wmem; // @[Core.scala 18:25]
  wire [31:0] reg_ex_wb_io_out_mem_addr; // @[Core.scala 18:25]
  wire [11:0] reg_ex_wb_io_out_aluop; // @[Core.scala 18:25]
  wire [6:0] reg_ex_wb_io_out_loadop; // @[Core.scala 18:25]
  wire [3:0] reg_ex_wb_io_out_storeop; // @[Core.scala 18:25]
  wire [3:0] reg_ex_wb_io_out_sysop; // @[Core.scala 18:25]
  wire  reg_ex_wb_io_out_bp_taken; // @[Core.scala 18:25]
  wire [31:0] reg_ex_wb_io_out_bp_targer; // @[Core.scala 18:25]
  wire  reg_ex_wb_io_stall; // @[Core.scala 18:25]
  wire  writeback_io_in_valid; // @[Core.scala 19:25]
  wire [31:0] writeback_io_in_pc; // @[Core.scala 19:25]
  wire [31:0] writeback_io_in_inst; // @[Core.scala 19:25]
  wire  writeback_io_in_wen; // @[Core.scala 19:25]
  wire [4:0] writeback_io_in_wdest; // @[Core.scala 19:25]
  wire [63:0] writeback_io_in_wdata; // @[Core.scala 19:25]
  wire [63:0] writeback_io_in_op1; // @[Core.scala 19:25]
  wire [31:0] writeback_io_in_mem_addr; // @[Core.scala 19:25]
  wire [6:0] writeback_io_in_loadop; // @[Core.scala 19:25]
  wire [3:0] writeback_io_in_storeop; // @[Core.scala 19:25]
  wire [3:0] writeback_io_in_sysop; // @[Core.scala 19:25]
  wire [31:0] writeback_io_pc; // @[Core.scala 19:25]
  wire [31:0] writeback_io_inst; // @[Core.scala 19:25]
  wire [63:0] writeback_io_op1; // @[Core.scala 19:25]
  wire [3:0] writeback_io_sysop; // @[Core.scala 19:25]
  wire [6:0] writeback_io_loadop; // @[Core.scala 19:25]
  wire [3:0] writeback_io_storeop; // @[Core.scala 19:25]
  wire [31:0] writeback_io_mem_addr; // @[Core.scala 19:25]
  wire  writeback_io_wen; // @[Core.scala 19:25]
  wire [4:0] writeback_io_wdest; // @[Core.scala 19:25]
  wire [63:0] writeback_io_wdata; // @[Core.scala 19:25]
  wire [4:0] writeback_io_wb_wdest; // @[Core.scala 19:25]
  wire [63:0] writeback_io_wb_result; // @[Core.scala 19:25]
  wire  writeback_io_exc; // @[Core.scala 19:25]
  wire  writeback_io_intr; // @[Core.scala 19:25]
  wire  writeback_io_ready_cmt; // @[Core.scala 19:25]
  wire  rf_clock; // @[Core.scala 20:18]
  wire  rf_reset; // @[Core.scala 20:18]
  wire [4:0] rf_io_rs1_addr; // @[Core.scala 20:18]
  wire [4:0] rf_io_rs2_addr; // @[Core.scala 20:18]
  wire [63:0] rf_io_rs1_data; // @[Core.scala 20:18]
  wire [63:0] rf_io_rs2_data; // @[Core.scala 20:18]
  wire  rf_io_wen; // @[Core.scala 20:18]
  wire [4:0] rf_io_wdest; // @[Core.scala 20:18]
  wire [63:0] rf_io_wdata; // @[Core.scala 20:18]
  wire [63:0] rf_rf_10; // @[Core.scala 20:18]
  wire  csr_clock; // @[Core.scala 21:19]
  wire  csr_reset; // @[Core.scala 21:19]
  wire [63:0] csr_io_in1; // @[Core.scala 21:19]
  wire [31:0] csr_io_pc; // @[Core.scala 21:19]
  wire [31:0] csr_io_inst; // @[Core.scala 21:19]
  wire [11:0] csr_io_raddr; // @[Core.scala 21:19]
  wire [3:0] csr_io_sysop; // @[Core.scala 21:19]
  wire  csr_io_exc; // @[Core.scala 21:19]
  wire [63:0] csr_io_csr_rdata; // @[Core.scala 21:19]
  wire [63:0] csr_io_mstatus; // @[Core.scala 21:19]
  wire [63:0] csr_io_mie; // @[Core.scala 21:19]
  wire [63:0] csr_io_mtvec; // @[Core.scala 21:19]
  wire [63:0] csr_io_mepc; // @[Core.scala 21:19]
  wire  clint_clock; // @[Core.scala 22:21]
  wire  clint_reset; // @[Core.scala 22:21]
  wire [63:0] clint_io_mstatus; // @[Core.scala 22:21]
  wire [63:0] clint_io_mie; // @[Core.scala 22:21]
  wire  clint_io_exc; // @[Core.scala 22:21]
  wire  clint_io_cmp_ren; // @[Core.scala 22:21]
  wire  clint_io_cmp_wen; // @[Core.scala 22:21]
  wire [63:0] clint_io_cmp_addr; // @[Core.scala 22:21]
  wire [63:0] clint_io_cmp_wdata; // @[Core.scala 22:21]
  wire [63:0] clint_io_cmp_rdata; // @[Core.scala 22:21]
  wire  clint_io_time_int; // @[Core.scala 22:21]
  wire  dt_ic_clock; // @[Core.scala 112:23]
  wire [7:0] dt_ic_coreid; // @[Core.scala 112:23]
  wire [7:0] dt_ic_index; // @[Core.scala 112:23]
  wire  dt_ic_valid; // @[Core.scala 112:23]
  wire [63:0] dt_ic_pc; // @[Core.scala 112:23]
  wire [31:0] dt_ic_instr; // @[Core.scala 112:23]
  wire [7:0] dt_ic_special; // @[Core.scala 112:23]
  wire  dt_ic_skip; // @[Core.scala 112:23]
  wire  dt_ic_isRVC; // @[Core.scala 112:23]
  wire  dt_ic_scFailed; // @[Core.scala 112:23]
  wire  dt_ic_wen; // @[Core.scala 112:23]
  wire [63:0] dt_ic_wdata; // @[Core.scala 112:23]
  wire [7:0] dt_ic_wdest; // @[Core.scala 112:23]
  wire  dt_ae_clock; // @[Core.scala 127:23]
  wire [7:0] dt_ae_coreid; // @[Core.scala 127:23]
  wire [31:0] dt_ae_intrNO; // @[Core.scala 127:23]
  wire [31:0] dt_ae_cause; // @[Core.scala 127:23]
  wire [63:0] dt_ae_exceptionPC; // @[Core.scala 127:23]
  wire [31:0] dt_ae_exceptionInst; // @[Core.scala 127:23]
  wire  dt_te_clock; // @[Core.scala 143:23]
  wire [7:0] dt_te_coreid; // @[Core.scala 143:23]
  wire  dt_te_valid; // @[Core.scala 143:23]
  wire [2:0] dt_te_code; // @[Core.scala 143:23]
  wire [63:0] dt_te_pc; // @[Core.scala 143:23]
  wire [63:0] dt_te_cycleCnt; // @[Core.scala 143:23]
  wire [63:0] dt_te_instrCnt; // @[Core.scala 143:23]
  wire  valid = writeback_io_ready_cmt & ~execution_io_busy; // @[Core.scala 86:40]
  wire [31:0] _inst_my_T = writeback_io_inst; // @[Core.scala 87:35]
  wire  inst_my = 32'h7b == _inst_my_T; // @[Core.scala 87:35]
  wire  _req_clint_T_5 = writeback_io_loadop != 7'h0 | writeback_io_storeop != 4'h0; // @[Core.scala 91:48]
  wire  req_clint = (writeback_io_mem_addr == 32'h2004000 | writeback_io_mem_addr == 32'h200bff8) & _req_clint_T_5; // @[Core.scala 90:103]
  reg  print_valid; // @[Core.scala 95:28]
  reg [63:0] print; // @[Core.scala 96:28]
  wire  _T = valid & inst_my; // @[Core.scala 97:15]
  reg  dt_ic_io_valid_REG; // @[Core.scala 116:33]
  reg [31:0] dt_ic_io_pc_REG; // @[Core.scala 117:33]
  reg [31:0] dt_ic_io_instr_REG; // @[Core.scala 118:33]
  reg  dt_ic_io_skip_REG; // @[Core.scala 120:33]
  reg  dt_ic_io_wen_REG; // @[Core.scala 123:33]
  reg [63:0] dt_ic_io_wdata_REG; // @[Core.scala 124:33]
  reg [4:0] dt_ic_io_wdest_REG; // @[Core.scala 125:33]
  reg [31:0] dt_ae_io_intrNO_REG; // @[Core.scala 130:37]
  reg [31:0] dt_ae_io_exceptionPC_REG; // @[Core.scala 132:37]
  reg [63:0] cycle_cnt; // @[Core.scala 134:28]
  reg [63:0] instr_cnt; // @[Core.scala 135:28]
  wire [63:0] _cycle_cnt_T_1 = cycle_cnt + 64'h1; // @[Core.scala 137:28]
  wire [63:0] _GEN_2 = {{63'd0}, valid}; // @[Core.scala 138:28]
  wire [63:0] _instr_cnt_T_1 = instr_cnt + _GEN_2; // @[Core.scala 138:28]
  wire [63:0] rf_a0_0 = rf_rf_10;
  InstFetch fetch ( // @[Core.scala 13:21]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_imem_inst_valid(fetch_io_imem_inst_valid),
    .io_imem_inst_ready(fetch_io_imem_inst_ready),
    .io_imem_inst_addr(fetch_io_imem_inst_addr),
    .io_imem_inst_read(fetch_io_imem_inst_read),
    .io_jmp_packet_valid(fetch_io_jmp_packet_valid),
    .io_jmp_packet_inst_pc(fetch_io_jmp_packet_inst_pc),
    .io_jmp_packet_jmp(fetch_io_jmp_packet_jmp),
    .io_jmp_packet_jmp_pc(fetch_io_jmp_packet_jmp_pc),
    .io_jmp_packet_mis(fetch_io_jmp_packet_mis),
    .io_stall(fetch_io_stall),
    .io_out_valid(fetch_io_out_valid),
    .io_out_pc(fetch_io_out_pc),
    .io_out_inst(fetch_io_out_inst),
    .io_out_bp_taken(fetch_io_out_bp_taken),
    .io_out_bp_targer(fetch_io_out_bp_targer)
  );
  PipelineReg reg_if_id ( // @[Core.scala 14:25]
    .clock(reg_if_id_clock),
    .reset(reg_if_id_reset),
    .io_in_valid(reg_if_id_io_in_valid),
    .io_in_pc(reg_if_id_io_in_pc),
    .io_in_inst(reg_if_id_io_in_inst),
    .io_in_wen(reg_if_id_io_in_wen),
    .io_in_wdest(reg_if_id_io_in_wdest),
    .io_in_wdata(reg_if_id_io_in_wdata),
    .io_in_op1(reg_if_id_io_in_op1),
    .io_in_op2(reg_if_id_io_in_op2),
    .io_in_typew(reg_if_id_io_in_typew),
    .io_in_wmem(reg_if_id_io_in_wmem),
    .io_in_mem_addr(reg_if_id_io_in_mem_addr),
    .io_in_aluop(reg_if_id_io_in_aluop),
    .io_in_loadop(reg_if_id_io_in_loadop),
    .io_in_storeop(reg_if_id_io_in_storeop),
    .io_in_sysop(reg_if_id_io_in_sysop),
    .io_in_bp_taken(reg_if_id_io_in_bp_taken),
    .io_in_bp_targer(reg_if_id_io_in_bp_targer),
    .io_out_valid(reg_if_id_io_out_valid),
    .io_out_pc(reg_if_id_io_out_pc),
    .io_out_inst(reg_if_id_io_out_inst),
    .io_out_wen(reg_if_id_io_out_wen),
    .io_out_wdest(reg_if_id_io_out_wdest),
    .io_out_wdata(reg_if_id_io_out_wdata),
    .io_out_op1(reg_if_id_io_out_op1),
    .io_out_op2(reg_if_id_io_out_op2),
    .io_out_typew(reg_if_id_io_out_typew),
    .io_out_wmem(reg_if_id_io_out_wmem),
    .io_out_mem_addr(reg_if_id_io_out_mem_addr),
    .io_out_aluop(reg_if_id_io_out_aluop),
    .io_out_loadop(reg_if_id_io_out_loadop),
    .io_out_storeop(reg_if_id_io_out_storeop),
    .io_out_sysop(reg_if_id_io_out_sysop),
    .io_out_bp_taken(reg_if_id_io_out_bp_taken),
    .io_out_bp_targer(reg_if_id_io_out_bp_targer),
    .io_stall(reg_if_id_io_stall)
  );
  Decode decode ( // @[Core.scala 15:22]
    .io_rs1_addr(decode_io_rs1_addr),
    .io_rs2_addr(decode_io_rs2_addr),
    .io_rs1_data(decode_io_rs1_data),
    .io_rs2_data(decode_io_rs2_data),
    .io_in_valid(decode_io_in_valid),
    .io_in_pc(decode_io_in_pc),
    .io_in_inst(decode_io_in_inst),
    .io_in_bp_taken(decode_io_in_bp_taken),
    .io_in_bp_targer(decode_io_in_bp_targer),
    .io_out_valid(decode_io_out_valid),
    .io_out_pc(decode_io_out_pc),
    .io_out_inst(decode_io_out_inst),
    .io_out_wen(decode_io_out_wen),
    .io_out_wdest(decode_io_out_wdest),
    .io_out_op1(decode_io_out_op1),
    .io_out_op2(decode_io_out_op2),
    .io_out_typew(decode_io_out_typew),
    .io_out_wmem(decode_io_out_wmem),
    .io_out_aluop(decode_io_out_aluop),
    .io_out_loadop(decode_io_out_loadop),
    .io_out_storeop(decode_io_out_storeop),
    .io_out_sysop(decode_io_out_sysop),
    .io_jmp_packet_valid(decode_io_jmp_packet_valid),
    .io_jmp_packet_inst_pc(decode_io_jmp_packet_inst_pc),
    .io_jmp_packet_jmp(decode_io_jmp_packet_jmp),
    .io_jmp_packet_jmp_pc(decode_io_jmp_packet_jmp_pc),
    .io_jmp_packet_mis(decode_io_jmp_packet_mis),
    .io_stall(decode_io_stall),
    .io_mtvec(decode_io_mtvec),
    .io_mepc(decode_io_mepc),
    .io_time_int(decode_io_time_int),
    .io_ex_wdest(decode_io_ex_wdest),
    .io_wb_wdest(decode_io_wb_wdest),
    .io_ex_result(decode_io_ex_result),
    .io_wb_result(decode_io_wb_result)
  );
  PipelineReg reg_id_ex ( // @[Core.scala 16:25]
    .clock(reg_id_ex_clock),
    .reset(reg_id_ex_reset),
    .io_in_valid(reg_id_ex_io_in_valid),
    .io_in_pc(reg_id_ex_io_in_pc),
    .io_in_inst(reg_id_ex_io_in_inst),
    .io_in_wen(reg_id_ex_io_in_wen),
    .io_in_wdest(reg_id_ex_io_in_wdest),
    .io_in_wdata(reg_id_ex_io_in_wdata),
    .io_in_op1(reg_id_ex_io_in_op1),
    .io_in_op2(reg_id_ex_io_in_op2),
    .io_in_typew(reg_id_ex_io_in_typew),
    .io_in_wmem(reg_id_ex_io_in_wmem),
    .io_in_mem_addr(reg_id_ex_io_in_mem_addr),
    .io_in_aluop(reg_id_ex_io_in_aluop),
    .io_in_loadop(reg_id_ex_io_in_loadop),
    .io_in_storeop(reg_id_ex_io_in_storeop),
    .io_in_sysop(reg_id_ex_io_in_sysop),
    .io_in_bp_taken(reg_id_ex_io_in_bp_taken),
    .io_in_bp_targer(reg_id_ex_io_in_bp_targer),
    .io_out_valid(reg_id_ex_io_out_valid),
    .io_out_pc(reg_id_ex_io_out_pc),
    .io_out_inst(reg_id_ex_io_out_inst),
    .io_out_wen(reg_id_ex_io_out_wen),
    .io_out_wdest(reg_id_ex_io_out_wdest),
    .io_out_wdata(reg_id_ex_io_out_wdata),
    .io_out_op1(reg_id_ex_io_out_op1),
    .io_out_op2(reg_id_ex_io_out_op2),
    .io_out_typew(reg_id_ex_io_out_typew),
    .io_out_wmem(reg_id_ex_io_out_wmem),
    .io_out_mem_addr(reg_id_ex_io_out_mem_addr),
    .io_out_aluop(reg_id_ex_io_out_aluop),
    .io_out_loadop(reg_id_ex_io_out_loadop),
    .io_out_storeop(reg_id_ex_io_out_storeop),
    .io_out_sysop(reg_id_ex_io_out_sysop),
    .io_out_bp_taken(reg_id_ex_io_out_bp_taken),
    .io_out_bp_targer(reg_id_ex_io_out_bp_targer),
    .io_stall(reg_id_ex_io_stall)
  );
  Execution execution ( // @[Core.scala 17:25]
    .clock(execution_clock),
    .reset(execution_reset),
    .io_in_valid(execution_io_in_valid),
    .io_in_pc(execution_io_in_pc),
    .io_in_inst(execution_io_in_inst),
    .io_in_wen(execution_io_in_wen),
    .io_in_wdest(execution_io_in_wdest),
    .io_in_op1(execution_io_in_op1),
    .io_in_op2(execution_io_in_op2),
    .io_in_typew(execution_io_in_typew),
    .io_in_wmem(execution_io_in_wmem),
    .io_in_aluop(execution_io_in_aluop),
    .io_in_loadop(execution_io_in_loadop),
    .io_in_storeop(execution_io_in_storeop),
    .io_in_sysop(execution_io_in_sysop),
    .io_out_valid(execution_io_out_valid),
    .io_out_pc(execution_io_out_pc),
    .io_out_inst(execution_io_out_inst),
    .io_out_wen(execution_io_out_wen),
    .io_out_wdest(execution_io_out_wdest),
    .io_out_wdata(execution_io_out_wdata),
    .io_out_op1(execution_io_out_op1),
    .io_out_op2(execution_io_out_op2),
    .io_out_typew(execution_io_out_typew),
    .io_out_wmem(execution_io_out_wmem),
    .io_out_mem_addr(execution_io_out_mem_addr),
    .io_out_aluop(execution_io_out_aluop),
    .io_out_loadop(execution_io_out_loadop),
    .io_out_storeop(execution_io_out_storeop),
    .io_out_sysop(execution_io_out_sysop),
    .io_busy(execution_io_busy),
    .io_csr_raddr(execution_io_csr_raddr),
    .io_csr_rdata(execution_io_csr_rdata),
    .io_dmem_data_valid(execution_io_dmem_data_valid),
    .io_dmem_data_ready(execution_io_dmem_data_ready),
    .io_dmem_data_req(execution_io_dmem_data_req),
    .io_dmem_data_addr(execution_io_dmem_data_addr),
    .io_dmem_data_size(execution_io_dmem_data_size),
    .io_dmem_data_strb(execution_io_dmem_data_strb),
    .io_dmem_data_read(execution_io_dmem_data_read),
    .io_dmem_data_write(execution_io_dmem_data_write),
    .io_cmp_ren(execution_io_cmp_ren),
    .io_cmp_wen(execution_io_cmp_wen),
    .io_cmp_addr(execution_io_cmp_addr),
    .io_cmp_wdata(execution_io_cmp_wdata),
    .io_cmp_rdata(execution_io_cmp_rdata),
    .io_ex_wdest(execution_io_ex_wdest),
    .io_ex_result(execution_io_ex_result)
  );
  PipelineReg reg_ex_wb ( // @[Core.scala 18:25]
    .clock(reg_ex_wb_clock),
    .reset(reg_ex_wb_reset),
    .io_in_valid(reg_ex_wb_io_in_valid),
    .io_in_pc(reg_ex_wb_io_in_pc),
    .io_in_inst(reg_ex_wb_io_in_inst),
    .io_in_wen(reg_ex_wb_io_in_wen),
    .io_in_wdest(reg_ex_wb_io_in_wdest),
    .io_in_wdata(reg_ex_wb_io_in_wdata),
    .io_in_op1(reg_ex_wb_io_in_op1),
    .io_in_op2(reg_ex_wb_io_in_op2),
    .io_in_typew(reg_ex_wb_io_in_typew),
    .io_in_wmem(reg_ex_wb_io_in_wmem),
    .io_in_mem_addr(reg_ex_wb_io_in_mem_addr),
    .io_in_aluop(reg_ex_wb_io_in_aluop),
    .io_in_loadop(reg_ex_wb_io_in_loadop),
    .io_in_storeop(reg_ex_wb_io_in_storeop),
    .io_in_sysop(reg_ex_wb_io_in_sysop),
    .io_in_bp_taken(reg_ex_wb_io_in_bp_taken),
    .io_in_bp_targer(reg_ex_wb_io_in_bp_targer),
    .io_out_valid(reg_ex_wb_io_out_valid),
    .io_out_pc(reg_ex_wb_io_out_pc),
    .io_out_inst(reg_ex_wb_io_out_inst),
    .io_out_wen(reg_ex_wb_io_out_wen),
    .io_out_wdest(reg_ex_wb_io_out_wdest),
    .io_out_wdata(reg_ex_wb_io_out_wdata),
    .io_out_op1(reg_ex_wb_io_out_op1),
    .io_out_op2(reg_ex_wb_io_out_op2),
    .io_out_typew(reg_ex_wb_io_out_typew),
    .io_out_wmem(reg_ex_wb_io_out_wmem),
    .io_out_mem_addr(reg_ex_wb_io_out_mem_addr),
    .io_out_aluop(reg_ex_wb_io_out_aluop),
    .io_out_loadop(reg_ex_wb_io_out_loadop),
    .io_out_storeop(reg_ex_wb_io_out_storeop),
    .io_out_sysop(reg_ex_wb_io_out_sysop),
    .io_out_bp_taken(reg_ex_wb_io_out_bp_taken),
    .io_out_bp_targer(reg_ex_wb_io_out_bp_targer),
    .io_stall(reg_ex_wb_io_stall)
  );
  WriteBack writeback ( // @[Core.scala 19:25]
    .io_in_valid(writeback_io_in_valid),
    .io_in_pc(writeback_io_in_pc),
    .io_in_inst(writeback_io_in_inst),
    .io_in_wen(writeback_io_in_wen),
    .io_in_wdest(writeback_io_in_wdest),
    .io_in_wdata(writeback_io_in_wdata),
    .io_in_op1(writeback_io_in_op1),
    .io_in_mem_addr(writeback_io_in_mem_addr),
    .io_in_loadop(writeback_io_in_loadop),
    .io_in_storeop(writeback_io_in_storeop),
    .io_in_sysop(writeback_io_in_sysop),
    .io_pc(writeback_io_pc),
    .io_inst(writeback_io_inst),
    .io_op1(writeback_io_op1),
    .io_sysop(writeback_io_sysop),
    .io_loadop(writeback_io_loadop),
    .io_storeop(writeback_io_storeop),
    .io_mem_addr(writeback_io_mem_addr),
    .io_wen(writeback_io_wen),
    .io_wdest(writeback_io_wdest),
    .io_wdata(writeback_io_wdata),
    .io_wb_wdest(writeback_io_wb_wdest),
    .io_wb_result(writeback_io_wb_result),
    .io_exc(writeback_io_exc),
    .io_intr(writeback_io_intr),
    .io_ready_cmt(writeback_io_ready_cmt)
  );
  RegFile rf ( // @[Core.scala 20:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_rs1_addr(rf_io_rs1_addr),
    .io_rs2_addr(rf_io_rs2_addr),
    .io_rs1_data(rf_io_rs1_data),
    .io_rs2_data(rf_io_rs2_data),
    .io_wen(rf_io_wen),
    .io_wdest(rf_io_wdest),
    .io_wdata(rf_io_wdata),
    .rf_10(rf_rf_10)
  );
  Csr csr ( // @[Core.scala 21:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in1(csr_io_in1),
    .io_pc(csr_io_pc),
    .io_inst(csr_io_inst),
    .io_raddr(csr_io_raddr),
    .io_sysop(csr_io_sysop),
    .io_exc(csr_io_exc),
    .io_csr_rdata(csr_io_csr_rdata),
    .io_mstatus(csr_io_mstatus),
    .io_mie(csr_io_mie),
    .io_mtvec(csr_io_mtvec),
    .io_mepc(csr_io_mepc)
  );
  Clint clint ( // @[Core.scala 22:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io_mstatus(clint_io_mstatus),
    .io_mie(clint_io_mie),
    .io_exc(clint_io_exc),
    .io_cmp_ren(clint_io_cmp_ren),
    .io_cmp_wen(clint_io_cmp_wen),
    .io_cmp_addr(clint_io_cmp_addr),
    .io_cmp_wdata(clint_io_cmp_wdata),
    .io_cmp_rdata(clint_io_cmp_rdata),
    .io_time_int(clint_io_time_int)
  );
  DifftestInstrCommit dt_ic ( // @[Core.scala 112:23]
    .clock(dt_ic_clock),
    .coreid(dt_ic_coreid),
    .index(dt_ic_index),
    .valid(dt_ic_valid),
    .pc(dt_ic_pc),
    .instr(dt_ic_instr),
    .special(dt_ic_special),
    .skip(dt_ic_skip),
    .isRVC(dt_ic_isRVC),
    .scFailed(dt_ic_scFailed),
    .wen(dt_ic_wen),
    .wdata(dt_ic_wdata),
    .wdest(dt_ic_wdest)
  );
  DifftestArchEvent dt_ae ( // @[Core.scala 127:23]
    .clock(dt_ae_clock),
    .coreid(dt_ae_coreid),
    .intrNO(dt_ae_intrNO),
    .cause(dt_ae_cause),
    .exceptionPC(dt_ae_exceptionPC),
    .exceptionInst(dt_ae_exceptionInst)
  );
  DifftestTrapEvent dt_te ( // @[Core.scala 143:23]
    .clock(dt_te_clock),
    .coreid(dt_te_coreid),
    .valid(dt_te_valid),
    .code(dt_te_code),
    .pc(dt_te_pc),
    .cycleCnt(dt_te_cycleCnt),
    .instrCnt(dt_te_instrCnt)
  );
  assign io_imem_inst_valid = fetch_io_imem_inst_valid; // @[Core.scala 27:27]
  assign io_imem_inst_addr = fetch_io_imem_inst_addr; // @[Core.scala 27:27]
  assign io_dmem_data_valid = execution_io_dmem_data_valid; // @[Core.scala 51:27]
  assign io_dmem_data_req = execution_io_dmem_data_req; // @[Core.scala 51:27]
  assign io_dmem_data_addr = execution_io_dmem_data_addr; // @[Core.scala 51:27]
  assign io_dmem_data_size = execution_io_dmem_data_size; // @[Core.scala 51:27]
  assign io_dmem_data_strb = execution_io_dmem_data_strb; // @[Core.scala 51:27]
  assign io_dmem_data_write = execution_io_dmem_data_write; // @[Core.scala 51:27]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_imem_inst_ready = io_imem_inst_ready; // @[Core.scala 27:27]
  assign fetch_io_imem_inst_read = io_imem_inst_read; // @[Core.scala 27:27]
  assign fetch_io_jmp_packet_valid = decode_io_jmp_packet_valid; // @[Core.scala 28:27]
  assign fetch_io_jmp_packet_inst_pc = decode_io_jmp_packet_inst_pc; // @[Core.scala 28:27]
  assign fetch_io_jmp_packet_jmp = decode_io_jmp_packet_jmp; // @[Core.scala 28:27]
  assign fetch_io_jmp_packet_jmp_pc = decode_io_jmp_packet_jmp_pc; // @[Core.scala 28:27]
  assign fetch_io_jmp_packet_mis = decode_io_jmp_packet_mis; // @[Core.scala 28:27]
  assign fetch_io_stall = execution_io_busy; // @[Core.scala 29:27]
  assign reg_if_id_clock = clock;
  assign reg_if_id_reset = reset;
  assign reg_if_id_io_in_valid = fetch_io_out_valid; // @[Core.scala 31:27]
  assign reg_if_id_io_in_pc = fetch_io_out_pc; // @[Core.scala 31:27]
  assign reg_if_id_io_in_inst = fetch_io_out_inst; // @[Core.scala 31:27]
  assign reg_if_id_io_in_wen = 1'h0; // @[Core.scala 31:27]
  assign reg_if_id_io_in_wdest = 5'h0; // @[Core.scala 31:27]
  assign reg_if_id_io_in_wdata = 64'h0; // @[Core.scala 31:27]
  assign reg_if_id_io_in_op1 = 64'h0; // @[Core.scala 31:27]
  assign reg_if_id_io_in_op2 = 64'h0; // @[Core.scala 31:27]
  assign reg_if_id_io_in_typew = 1'h0; // @[Core.scala 31:27]
  assign reg_if_id_io_in_wmem = 64'h0; // @[Core.scala 31:27]
  assign reg_if_id_io_in_mem_addr = 32'h0; // @[Core.scala 31:27]
  assign reg_if_id_io_in_aluop = 12'h0; // @[Core.scala 31:27]
  assign reg_if_id_io_in_loadop = 7'h0; // @[Core.scala 31:27]
  assign reg_if_id_io_in_storeop = 4'h0; // @[Core.scala 31:27]
  assign reg_if_id_io_in_sysop = 4'h0; // @[Core.scala 31:27]
  assign reg_if_id_io_in_bp_taken = fetch_io_out_bp_taken; // @[Core.scala 31:27]
  assign reg_if_id_io_in_bp_targer = fetch_io_out_bp_targer; // @[Core.scala 31:27]
  assign reg_if_id_io_stall = execution_io_busy; // @[Core.scala 32:27]
  assign decode_io_rs1_data = rf_io_rs1_data; // @[Core.scala 36:27]
  assign decode_io_rs2_data = rf_io_rs2_data; // @[Core.scala 37:27]
  assign decode_io_in_valid = reg_if_id_io_out_valid; // @[Core.scala 35:27]
  assign decode_io_in_pc = reg_if_id_io_out_pc; // @[Core.scala 35:27]
  assign decode_io_in_inst = reg_if_id_io_out_inst; // @[Core.scala 35:27]
  assign decode_io_in_bp_taken = reg_if_id_io_out_bp_taken; // @[Core.scala 35:27]
  assign decode_io_in_bp_targer = reg_if_id_io_out_bp_targer; // @[Core.scala 35:27]
  assign decode_io_stall = execution_io_busy; // @[Core.scala 38:27]
  assign decode_io_mtvec = csr_io_mtvec; // @[Core.scala 43:27]
  assign decode_io_mepc = csr_io_mepc; // @[Core.scala 44:27]
  assign decode_io_time_int = clint_io_time_int; // @[Core.scala 45:27]
  assign decode_io_ex_wdest = execution_io_ex_wdest; // @[Core.scala 39:27]
  assign decode_io_wb_wdest = writeback_io_wb_wdest; // @[Core.scala 41:27]
  assign decode_io_ex_result = execution_io_ex_result; // @[Core.scala 40:27]
  assign decode_io_wb_result = writeback_io_wb_result; // @[Core.scala 42:27]
  assign reg_id_ex_clock = clock;
  assign reg_id_ex_reset = reset;
  assign reg_id_ex_io_in_valid = decode_io_out_valid; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_pc = decode_io_out_pc; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_inst = decode_io_out_inst; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_wen = decode_io_out_wen; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_wdest = decode_io_out_wdest; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_wdata = 64'h0; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_op1 = decode_io_out_op1; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_op2 = decode_io_out_op2; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_typew = decode_io_out_typew; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_wmem = decode_io_out_wmem; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_mem_addr = 32'h0; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_aluop = decode_io_out_aluop; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_loadop = decode_io_out_loadop; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_storeop = decode_io_out_storeop; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_sysop = decode_io_out_sysop; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_bp_taken = 1'h0; // @[Core.scala 47:27]
  assign reg_id_ex_io_in_bp_targer = 32'h0; // @[Core.scala 47:27]
  assign reg_id_ex_io_stall = execution_io_busy; // @[Core.scala 48:27]
  assign execution_clock = clock;
  assign execution_reset = reset;
  assign execution_io_in_valid = reg_id_ex_io_out_valid; // @[Core.scala 52:27]
  assign execution_io_in_pc = reg_id_ex_io_out_pc; // @[Core.scala 52:27]
  assign execution_io_in_inst = reg_id_ex_io_out_inst; // @[Core.scala 52:27]
  assign execution_io_in_wen = reg_id_ex_io_out_wen; // @[Core.scala 52:27]
  assign execution_io_in_wdest = reg_id_ex_io_out_wdest; // @[Core.scala 52:27]
  assign execution_io_in_op1 = reg_id_ex_io_out_op1; // @[Core.scala 52:27]
  assign execution_io_in_op2 = reg_id_ex_io_out_op2; // @[Core.scala 52:27]
  assign execution_io_in_typew = reg_id_ex_io_out_typew; // @[Core.scala 52:27]
  assign execution_io_in_wmem = reg_id_ex_io_out_wmem; // @[Core.scala 52:27]
  assign execution_io_in_aluop = reg_id_ex_io_out_aluop; // @[Core.scala 52:27]
  assign execution_io_in_loadop = reg_id_ex_io_out_loadop; // @[Core.scala 52:27]
  assign execution_io_in_storeop = reg_id_ex_io_out_storeop; // @[Core.scala 52:27]
  assign execution_io_in_sysop = reg_id_ex_io_out_sysop; // @[Core.scala 52:27]
  assign execution_io_csr_rdata = csr_io_csr_rdata; // @[Core.scala 53:27]
  assign execution_io_dmem_data_ready = io_dmem_data_ready; // @[Core.scala 51:27]
  assign execution_io_dmem_data_read = io_dmem_data_read; // @[Core.scala 51:27]
  assign execution_io_cmp_rdata = clint_io_cmp_rdata; // @[Core.scala 54:27]
  assign reg_ex_wb_clock = clock;
  assign reg_ex_wb_reset = reset;
  assign reg_ex_wb_io_in_valid = execution_io_out_valid; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_pc = execution_io_out_pc; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_inst = execution_io_out_inst; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_wen = execution_io_out_wen; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_wdest = execution_io_out_wdest; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_wdata = execution_io_out_wdata; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_op1 = execution_io_out_op1; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_op2 = execution_io_out_op2; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_typew = execution_io_out_typew; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_wmem = execution_io_out_wmem; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_mem_addr = execution_io_out_mem_addr; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_aluop = execution_io_out_aluop; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_loadop = execution_io_out_loadop; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_storeop = execution_io_out_storeop; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_sysop = execution_io_out_sysop; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_bp_taken = 1'h0; // @[Core.scala 56:27]
  assign reg_ex_wb_io_in_bp_targer = 32'h0; // @[Core.scala 56:27]
  assign reg_ex_wb_io_stall = execution_io_busy; // @[Core.scala 57:27]
  assign writeback_io_in_valid = reg_ex_wb_io_out_valid; // @[Core.scala 60:27]
  assign writeback_io_in_pc = reg_ex_wb_io_out_pc; // @[Core.scala 60:27]
  assign writeback_io_in_inst = reg_ex_wb_io_out_inst; // @[Core.scala 60:27]
  assign writeback_io_in_wen = reg_ex_wb_io_out_wen; // @[Core.scala 60:27]
  assign writeback_io_in_wdest = reg_ex_wb_io_out_wdest; // @[Core.scala 60:27]
  assign writeback_io_in_wdata = reg_ex_wb_io_out_wdata; // @[Core.scala 60:27]
  assign writeback_io_in_op1 = reg_ex_wb_io_out_op1; // @[Core.scala 60:27]
  assign writeback_io_in_mem_addr = reg_ex_wb_io_out_mem_addr; // @[Core.scala 60:27]
  assign writeback_io_in_loadop = reg_ex_wb_io_out_loadop; // @[Core.scala 60:27]
  assign writeback_io_in_storeop = reg_ex_wb_io_out_storeop; // @[Core.scala 60:27]
  assign writeback_io_in_sysop = reg_ex_wb_io_out_sysop; // @[Core.scala 60:27]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_rs1_addr = decode_io_rs1_addr; // @[Core.scala 62:27]
  assign rf_io_rs2_addr = decode_io_rs2_addr; // @[Core.scala 63:27]
  assign rf_io_wen = writeback_io_wen; // @[Core.scala 64:27]
  assign rf_io_wdest = writeback_io_wdest; // @[Core.scala 65:27]
  assign rf_io_wdata = writeback_io_wdata; // @[Core.scala 66:27]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in1 = writeback_io_op1; // @[Core.scala 68:27]
  assign csr_io_pc = writeback_io_pc; // @[Core.scala 72:27]
  assign csr_io_inst = writeback_io_inst; // @[Core.scala 71:27]
  assign csr_io_raddr = execution_io_csr_raddr; // @[Core.scala 70:27]
  assign csr_io_sysop = writeback_io_sysop; // @[Core.scala 69:27]
  assign csr_io_exc = writeback_io_exc; // @[Core.scala 73:27]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io_mstatus = csr_io_mstatus; // @[Core.scala 75:27]
  assign clint_io_mie = csr_io_mie; // @[Core.scala 76:27]
  assign clint_io_exc = writeback_io_exc; // @[Core.scala 77:27]
  assign clint_io_cmp_ren = execution_io_cmp_ren; // @[Core.scala 78:27]
  assign clint_io_cmp_wen = execution_io_cmp_wen; // @[Core.scala 79:27]
  assign clint_io_cmp_addr = execution_io_cmp_addr; // @[Core.scala 80:27]
  assign clint_io_cmp_wdata = execution_io_cmp_wdata; // @[Core.scala 81:27]
  assign dt_ic_clock = clock; // @[Core.scala 113:23]
  assign dt_ic_coreid = 8'h0; // @[Core.scala 114:23]
  assign dt_ic_index = 8'h0; // @[Core.scala 115:23]
  assign dt_ic_valid = dt_ic_io_valid_REG; // @[Core.scala 116:23]
  assign dt_ic_pc = {{32'd0}, dt_ic_io_pc_REG}; // @[Core.scala 117:23]
  assign dt_ic_instr = dt_ic_io_instr_REG; // @[Core.scala 118:23]
  assign dt_ic_special = 8'h0; // @[Core.scala 119:23]
  assign dt_ic_skip = dt_ic_io_skip_REG; // @[Core.scala 120:23]
  assign dt_ic_isRVC = 1'h0; // @[Core.scala 121:23]
  assign dt_ic_scFailed = 1'h0; // @[Core.scala 122:23]
  assign dt_ic_wen = dt_ic_io_wen_REG; // @[Core.scala 123:23]
  assign dt_ic_wdata = dt_ic_io_wdata_REG; // @[Core.scala 124:23]
  assign dt_ic_wdest = {{3'd0}, dt_ic_io_wdest_REG}; // @[Core.scala 125:23]
  assign dt_ae_clock = clock; // @[Core.scala 128:27]
  assign dt_ae_coreid = 8'h0; // @[Core.scala 129:27]
  assign dt_ae_intrNO = dt_ae_io_intrNO_REG; // @[Core.scala 130:27]
  assign dt_ae_cause = 32'h0; // @[Core.scala 131:27]
  assign dt_ae_exceptionPC = {{32'd0}, dt_ae_io_exceptionPC_REG}; // @[Core.scala 132:27]
  assign dt_ae_exceptionInst = 32'h0;
  assign dt_te_clock = clock; // @[Core.scala 144:23]
  assign dt_te_coreid = 8'h0; // @[Core.scala 145:23]
  assign dt_te_valid = writeback_io_inst == 32'h6b; // @[Core.scala 146:45]
  assign dt_te_code = rf_a0_0[2:0]; // @[Core.scala 147:31]
  assign dt_te_pc = {{32'd0}, writeback_io_pc}; // @[Core.scala 148:23]
  assign dt_te_cycleCnt = cycle_cnt; // @[Core.scala 149:23]
  assign dt_te_instrCnt = instr_cnt; // @[Core.scala 150:23]
  always @(posedge clock) begin
    if (reset) begin // @[Core.scala 95:28]
      print_valid <= 1'h0; // @[Core.scala 95:28]
    end else begin
      print_valid <= _T;
    end
    if (reset) begin // @[Core.scala 96:28]
      print <= 64'h0; // @[Core.scala 96:28]
    end else if (valid & inst_my) begin // @[Core.scala 97:27]
      print <= writeback_io_op1; // @[Core.scala 99:11]
    end
    dt_ic_io_valid_REG <= writeback_io_ready_cmt & ~execution_io_busy; // @[Core.scala 86:40]
    dt_ic_io_pc_REG <= writeback_io_pc; // @[Core.scala 117:33]
    dt_ic_io_instr_REG <= writeback_io_inst; // @[Core.scala 118:33]
    dt_ic_io_skip_REG <= inst_my | writeback_io_inst[31:20] == 12'hb00 & writeback_io_sysop != 4'h0 | req_clint; // @[Core.scala 93:102]
    dt_ic_io_wen_REG <= writeback_io_wen; // @[Core.scala 123:33]
    dt_ic_io_wdata_REG <= writeback_io_wdata; // @[Core.scala 124:33]
    dt_ic_io_wdest_REG <= writeback_io_wdest; // @[Core.scala 125:33]
    if (writeback_io_intr) begin // @[Core.scala 108:20]
      dt_ae_io_intrNO_REG <= 32'h7;
    end else begin
      dt_ae_io_intrNO_REG <= 32'h0;
    end
    if (writeback_io_intr) begin // @[Core.scala 109:24]
      dt_ae_io_exceptionPC_REG <= writeback_io_pc;
    end else begin
      dt_ae_io_exceptionPC_REG <= 32'h0;
    end
    if (reset) begin // @[Core.scala 134:28]
      cycle_cnt <= 64'h0; // @[Core.scala 134:28]
    end else begin
      cycle_cnt <= _cycle_cnt_T_1; // @[Core.scala 137:15]
    end
    if (reset) begin // @[Core.scala 135:28]
      instr_cnt <= 64'h0; // @[Core.scala 135:28]
    end else begin
      instr_cnt <= _instr_cnt_T_1; // @[Core.scala 138:15]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (print_valid & ~reset) begin
          $fwrite(32'h80000002,"%c",print); // @[Core.scala 104:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  print_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  print = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  dt_ic_io_valid_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  dt_ic_io_pc_REG = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  dt_ic_io_instr_REG = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  dt_ic_io_skip_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dt_ic_io_wen_REG = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  dt_ic_io_wdata_REG = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  dt_ic_io_wdest_REG = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  dt_ae_io_intrNO_REG = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  dt_ae_io_exceptionPC_REG = _RAND_10[31:0];
  _RAND_11 = {2{`RANDOM}};
  cycle_cnt = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  instr_cnt = _RAND_12[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Icache(
  input          clock,
  input          reset,
  input          io_imem_inst_valid,
  output         io_imem_inst_ready,
  input  [31:0]  io_imem_inst_addr,
  output [31:0]  io_imem_inst_read,
  output         io_out_inst_valid,
  input          io_out_inst_ready,
  output [31:0]  io_out_inst_addr,
  input  [127:0] io_out_inst_read
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [127:0] _RAND_516;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] req_Q; // @[Icache.scala 114:19]
  wire  req_CLK; // @[Icache.scala 114:19]
  wire  req_CEN; // @[Icache.scala 114:19]
  wire  req_WEN; // @[Icache.scala 114:19]
  wire [7:0] req_A; // @[Icache.scala 114:19]
  wire [127:0] req_D; // @[Icache.scala 114:19]
  reg [19:0] tag_0; // @[Icache.scala 16:24]
  reg [19:0] tag_1; // @[Icache.scala 16:24]
  reg [19:0] tag_2; // @[Icache.scala 16:24]
  reg [19:0] tag_3; // @[Icache.scala 16:24]
  reg [19:0] tag_4; // @[Icache.scala 16:24]
  reg [19:0] tag_5; // @[Icache.scala 16:24]
  reg [19:0] tag_6; // @[Icache.scala 16:24]
  reg [19:0] tag_7; // @[Icache.scala 16:24]
  reg [19:0] tag_8; // @[Icache.scala 16:24]
  reg [19:0] tag_9; // @[Icache.scala 16:24]
  reg [19:0] tag_10; // @[Icache.scala 16:24]
  reg [19:0] tag_11; // @[Icache.scala 16:24]
  reg [19:0] tag_12; // @[Icache.scala 16:24]
  reg [19:0] tag_13; // @[Icache.scala 16:24]
  reg [19:0] tag_14; // @[Icache.scala 16:24]
  reg [19:0] tag_15; // @[Icache.scala 16:24]
  reg [19:0] tag_16; // @[Icache.scala 16:24]
  reg [19:0] tag_17; // @[Icache.scala 16:24]
  reg [19:0] tag_18; // @[Icache.scala 16:24]
  reg [19:0] tag_19; // @[Icache.scala 16:24]
  reg [19:0] tag_20; // @[Icache.scala 16:24]
  reg [19:0] tag_21; // @[Icache.scala 16:24]
  reg [19:0] tag_22; // @[Icache.scala 16:24]
  reg [19:0] tag_23; // @[Icache.scala 16:24]
  reg [19:0] tag_24; // @[Icache.scala 16:24]
  reg [19:0] tag_25; // @[Icache.scala 16:24]
  reg [19:0] tag_26; // @[Icache.scala 16:24]
  reg [19:0] tag_27; // @[Icache.scala 16:24]
  reg [19:0] tag_28; // @[Icache.scala 16:24]
  reg [19:0] tag_29; // @[Icache.scala 16:24]
  reg [19:0] tag_30; // @[Icache.scala 16:24]
  reg [19:0] tag_31; // @[Icache.scala 16:24]
  reg [19:0] tag_32; // @[Icache.scala 16:24]
  reg [19:0] tag_33; // @[Icache.scala 16:24]
  reg [19:0] tag_34; // @[Icache.scala 16:24]
  reg [19:0] tag_35; // @[Icache.scala 16:24]
  reg [19:0] tag_36; // @[Icache.scala 16:24]
  reg [19:0] tag_37; // @[Icache.scala 16:24]
  reg [19:0] tag_38; // @[Icache.scala 16:24]
  reg [19:0] tag_39; // @[Icache.scala 16:24]
  reg [19:0] tag_40; // @[Icache.scala 16:24]
  reg [19:0] tag_41; // @[Icache.scala 16:24]
  reg [19:0] tag_42; // @[Icache.scala 16:24]
  reg [19:0] tag_43; // @[Icache.scala 16:24]
  reg [19:0] tag_44; // @[Icache.scala 16:24]
  reg [19:0] tag_45; // @[Icache.scala 16:24]
  reg [19:0] tag_46; // @[Icache.scala 16:24]
  reg [19:0] tag_47; // @[Icache.scala 16:24]
  reg [19:0] tag_48; // @[Icache.scala 16:24]
  reg [19:0] tag_49; // @[Icache.scala 16:24]
  reg [19:0] tag_50; // @[Icache.scala 16:24]
  reg [19:0] tag_51; // @[Icache.scala 16:24]
  reg [19:0] tag_52; // @[Icache.scala 16:24]
  reg [19:0] tag_53; // @[Icache.scala 16:24]
  reg [19:0] tag_54; // @[Icache.scala 16:24]
  reg [19:0] tag_55; // @[Icache.scala 16:24]
  reg [19:0] tag_56; // @[Icache.scala 16:24]
  reg [19:0] tag_57; // @[Icache.scala 16:24]
  reg [19:0] tag_58; // @[Icache.scala 16:24]
  reg [19:0] tag_59; // @[Icache.scala 16:24]
  reg [19:0] tag_60; // @[Icache.scala 16:24]
  reg [19:0] tag_61; // @[Icache.scala 16:24]
  reg [19:0] tag_62; // @[Icache.scala 16:24]
  reg [19:0] tag_63; // @[Icache.scala 16:24]
  reg [19:0] tag_64; // @[Icache.scala 16:24]
  reg [19:0] tag_65; // @[Icache.scala 16:24]
  reg [19:0] tag_66; // @[Icache.scala 16:24]
  reg [19:0] tag_67; // @[Icache.scala 16:24]
  reg [19:0] tag_68; // @[Icache.scala 16:24]
  reg [19:0] tag_69; // @[Icache.scala 16:24]
  reg [19:0] tag_70; // @[Icache.scala 16:24]
  reg [19:0] tag_71; // @[Icache.scala 16:24]
  reg [19:0] tag_72; // @[Icache.scala 16:24]
  reg [19:0] tag_73; // @[Icache.scala 16:24]
  reg [19:0] tag_74; // @[Icache.scala 16:24]
  reg [19:0] tag_75; // @[Icache.scala 16:24]
  reg [19:0] tag_76; // @[Icache.scala 16:24]
  reg [19:0] tag_77; // @[Icache.scala 16:24]
  reg [19:0] tag_78; // @[Icache.scala 16:24]
  reg [19:0] tag_79; // @[Icache.scala 16:24]
  reg [19:0] tag_80; // @[Icache.scala 16:24]
  reg [19:0] tag_81; // @[Icache.scala 16:24]
  reg [19:0] tag_82; // @[Icache.scala 16:24]
  reg [19:0] tag_83; // @[Icache.scala 16:24]
  reg [19:0] tag_84; // @[Icache.scala 16:24]
  reg [19:0] tag_85; // @[Icache.scala 16:24]
  reg [19:0] tag_86; // @[Icache.scala 16:24]
  reg [19:0] tag_87; // @[Icache.scala 16:24]
  reg [19:0] tag_88; // @[Icache.scala 16:24]
  reg [19:0] tag_89; // @[Icache.scala 16:24]
  reg [19:0] tag_90; // @[Icache.scala 16:24]
  reg [19:0] tag_91; // @[Icache.scala 16:24]
  reg [19:0] tag_92; // @[Icache.scala 16:24]
  reg [19:0] tag_93; // @[Icache.scala 16:24]
  reg [19:0] tag_94; // @[Icache.scala 16:24]
  reg [19:0] tag_95; // @[Icache.scala 16:24]
  reg [19:0] tag_96; // @[Icache.scala 16:24]
  reg [19:0] tag_97; // @[Icache.scala 16:24]
  reg [19:0] tag_98; // @[Icache.scala 16:24]
  reg [19:0] tag_99; // @[Icache.scala 16:24]
  reg [19:0] tag_100; // @[Icache.scala 16:24]
  reg [19:0] tag_101; // @[Icache.scala 16:24]
  reg [19:0] tag_102; // @[Icache.scala 16:24]
  reg [19:0] tag_103; // @[Icache.scala 16:24]
  reg [19:0] tag_104; // @[Icache.scala 16:24]
  reg [19:0] tag_105; // @[Icache.scala 16:24]
  reg [19:0] tag_106; // @[Icache.scala 16:24]
  reg [19:0] tag_107; // @[Icache.scala 16:24]
  reg [19:0] tag_108; // @[Icache.scala 16:24]
  reg [19:0] tag_109; // @[Icache.scala 16:24]
  reg [19:0] tag_110; // @[Icache.scala 16:24]
  reg [19:0] tag_111; // @[Icache.scala 16:24]
  reg [19:0] tag_112; // @[Icache.scala 16:24]
  reg [19:0] tag_113; // @[Icache.scala 16:24]
  reg [19:0] tag_114; // @[Icache.scala 16:24]
  reg [19:0] tag_115; // @[Icache.scala 16:24]
  reg [19:0] tag_116; // @[Icache.scala 16:24]
  reg [19:0] tag_117; // @[Icache.scala 16:24]
  reg [19:0] tag_118; // @[Icache.scala 16:24]
  reg [19:0] tag_119; // @[Icache.scala 16:24]
  reg [19:0] tag_120; // @[Icache.scala 16:24]
  reg [19:0] tag_121; // @[Icache.scala 16:24]
  reg [19:0] tag_122; // @[Icache.scala 16:24]
  reg [19:0] tag_123; // @[Icache.scala 16:24]
  reg [19:0] tag_124; // @[Icache.scala 16:24]
  reg [19:0] tag_125; // @[Icache.scala 16:24]
  reg [19:0] tag_126; // @[Icache.scala 16:24]
  reg [19:0] tag_127; // @[Icache.scala 16:24]
  reg [19:0] tag_128; // @[Icache.scala 16:24]
  reg [19:0] tag_129; // @[Icache.scala 16:24]
  reg [19:0] tag_130; // @[Icache.scala 16:24]
  reg [19:0] tag_131; // @[Icache.scala 16:24]
  reg [19:0] tag_132; // @[Icache.scala 16:24]
  reg [19:0] tag_133; // @[Icache.scala 16:24]
  reg [19:0] tag_134; // @[Icache.scala 16:24]
  reg [19:0] tag_135; // @[Icache.scala 16:24]
  reg [19:0] tag_136; // @[Icache.scala 16:24]
  reg [19:0] tag_137; // @[Icache.scala 16:24]
  reg [19:0] tag_138; // @[Icache.scala 16:24]
  reg [19:0] tag_139; // @[Icache.scala 16:24]
  reg [19:0] tag_140; // @[Icache.scala 16:24]
  reg [19:0] tag_141; // @[Icache.scala 16:24]
  reg [19:0] tag_142; // @[Icache.scala 16:24]
  reg [19:0] tag_143; // @[Icache.scala 16:24]
  reg [19:0] tag_144; // @[Icache.scala 16:24]
  reg [19:0] tag_145; // @[Icache.scala 16:24]
  reg [19:0] tag_146; // @[Icache.scala 16:24]
  reg [19:0] tag_147; // @[Icache.scala 16:24]
  reg [19:0] tag_148; // @[Icache.scala 16:24]
  reg [19:0] tag_149; // @[Icache.scala 16:24]
  reg [19:0] tag_150; // @[Icache.scala 16:24]
  reg [19:0] tag_151; // @[Icache.scala 16:24]
  reg [19:0] tag_152; // @[Icache.scala 16:24]
  reg [19:0] tag_153; // @[Icache.scala 16:24]
  reg [19:0] tag_154; // @[Icache.scala 16:24]
  reg [19:0] tag_155; // @[Icache.scala 16:24]
  reg [19:0] tag_156; // @[Icache.scala 16:24]
  reg [19:0] tag_157; // @[Icache.scala 16:24]
  reg [19:0] tag_158; // @[Icache.scala 16:24]
  reg [19:0] tag_159; // @[Icache.scala 16:24]
  reg [19:0] tag_160; // @[Icache.scala 16:24]
  reg [19:0] tag_161; // @[Icache.scala 16:24]
  reg [19:0] tag_162; // @[Icache.scala 16:24]
  reg [19:0] tag_163; // @[Icache.scala 16:24]
  reg [19:0] tag_164; // @[Icache.scala 16:24]
  reg [19:0] tag_165; // @[Icache.scala 16:24]
  reg [19:0] tag_166; // @[Icache.scala 16:24]
  reg [19:0] tag_167; // @[Icache.scala 16:24]
  reg [19:0] tag_168; // @[Icache.scala 16:24]
  reg [19:0] tag_169; // @[Icache.scala 16:24]
  reg [19:0] tag_170; // @[Icache.scala 16:24]
  reg [19:0] tag_171; // @[Icache.scala 16:24]
  reg [19:0] tag_172; // @[Icache.scala 16:24]
  reg [19:0] tag_173; // @[Icache.scala 16:24]
  reg [19:0] tag_174; // @[Icache.scala 16:24]
  reg [19:0] tag_175; // @[Icache.scala 16:24]
  reg [19:0] tag_176; // @[Icache.scala 16:24]
  reg [19:0] tag_177; // @[Icache.scala 16:24]
  reg [19:0] tag_178; // @[Icache.scala 16:24]
  reg [19:0] tag_179; // @[Icache.scala 16:24]
  reg [19:0] tag_180; // @[Icache.scala 16:24]
  reg [19:0] tag_181; // @[Icache.scala 16:24]
  reg [19:0] tag_182; // @[Icache.scala 16:24]
  reg [19:0] tag_183; // @[Icache.scala 16:24]
  reg [19:0] tag_184; // @[Icache.scala 16:24]
  reg [19:0] tag_185; // @[Icache.scala 16:24]
  reg [19:0] tag_186; // @[Icache.scala 16:24]
  reg [19:0] tag_187; // @[Icache.scala 16:24]
  reg [19:0] tag_188; // @[Icache.scala 16:24]
  reg [19:0] tag_189; // @[Icache.scala 16:24]
  reg [19:0] tag_190; // @[Icache.scala 16:24]
  reg [19:0] tag_191; // @[Icache.scala 16:24]
  reg [19:0] tag_192; // @[Icache.scala 16:24]
  reg [19:0] tag_193; // @[Icache.scala 16:24]
  reg [19:0] tag_194; // @[Icache.scala 16:24]
  reg [19:0] tag_195; // @[Icache.scala 16:24]
  reg [19:0] tag_196; // @[Icache.scala 16:24]
  reg [19:0] tag_197; // @[Icache.scala 16:24]
  reg [19:0] tag_198; // @[Icache.scala 16:24]
  reg [19:0] tag_199; // @[Icache.scala 16:24]
  reg [19:0] tag_200; // @[Icache.scala 16:24]
  reg [19:0] tag_201; // @[Icache.scala 16:24]
  reg [19:0] tag_202; // @[Icache.scala 16:24]
  reg [19:0] tag_203; // @[Icache.scala 16:24]
  reg [19:0] tag_204; // @[Icache.scala 16:24]
  reg [19:0] tag_205; // @[Icache.scala 16:24]
  reg [19:0] tag_206; // @[Icache.scala 16:24]
  reg [19:0] tag_207; // @[Icache.scala 16:24]
  reg [19:0] tag_208; // @[Icache.scala 16:24]
  reg [19:0] tag_209; // @[Icache.scala 16:24]
  reg [19:0] tag_210; // @[Icache.scala 16:24]
  reg [19:0] tag_211; // @[Icache.scala 16:24]
  reg [19:0] tag_212; // @[Icache.scala 16:24]
  reg [19:0] tag_213; // @[Icache.scala 16:24]
  reg [19:0] tag_214; // @[Icache.scala 16:24]
  reg [19:0] tag_215; // @[Icache.scala 16:24]
  reg [19:0] tag_216; // @[Icache.scala 16:24]
  reg [19:0] tag_217; // @[Icache.scala 16:24]
  reg [19:0] tag_218; // @[Icache.scala 16:24]
  reg [19:0] tag_219; // @[Icache.scala 16:24]
  reg [19:0] tag_220; // @[Icache.scala 16:24]
  reg [19:0] tag_221; // @[Icache.scala 16:24]
  reg [19:0] tag_222; // @[Icache.scala 16:24]
  reg [19:0] tag_223; // @[Icache.scala 16:24]
  reg [19:0] tag_224; // @[Icache.scala 16:24]
  reg [19:0] tag_225; // @[Icache.scala 16:24]
  reg [19:0] tag_226; // @[Icache.scala 16:24]
  reg [19:0] tag_227; // @[Icache.scala 16:24]
  reg [19:0] tag_228; // @[Icache.scala 16:24]
  reg [19:0] tag_229; // @[Icache.scala 16:24]
  reg [19:0] tag_230; // @[Icache.scala 16:24]
  reg [19:0] tag_231; // @[Icache.scala 16:24]
  reg [19:0] tag_232; // @[Icache.scala 16:24]
  reg [19:0] tag_233; // @[Icache.scala 16:24]
  reg [19:0] tag_234; // @[Icache.scala 16:24]
  reg [19:0] tag_235; // @[Icache.scala 16:24]
  reg [19:0] tag_236; // @[Icache.scala 16:24]
  reg [19:0] tag_237; // @[Icache.scala 16:24]
  reg [19:0] tag_238; // @[Icache.scala 16:24]
  reg [19:0] tag_239; // @[Icache.scala 16:24]
  reg [19:0] tag_240; // @[Icache.scala 16:24]
  reg [19:0] tag_241; // @[Icache.scala 16:24]
  reg [19:0] tag_242; // @[Icache.scala 16:24]
  reg [19:0] tag_243; // @[Icache.scala 16:24]
  reg [19:0] tag_244; // @[Icache.scala 16:24]
  reg [19:0] tag_245; // @[Icache.scala 16:24]
  reg [19:0] tag_246; // @[Icache.scala 16:24]
  reg [19:0] tag_247; // @[Icache.scala 16:24]
  reg [19:0] tag_248; // @[Icache.scala 16:24]
  reg [19:0] tag_249; // @[Icache.scala 16:24]
  reg [19:0] tag_250; // @[Icache.scala 16:24]
  reg [19:0] tag_251; // @[Icache.scala 16:24]
  reg [19:0] tag_252; // @[Icache.scala 16:24]
  reg [19:0] tag_253; // @[Icache.scala 16:24]
  reg [19:0] tag_254; // @[Icache.scala 16:24]
  reg [19:0] tag_255; // @[Icache.scala 16:24]
  reg  valid_0; // @[Icache.scala 17:24]
  reg  valid_1; // @[Icache.scala 17:24]
  reg  valid_2; // @[Icache.scala 17:24]
  reg  valid_3; // @[Icache.scala 17:24]
  reg  valid_4; // @[Icache.scala 17:24]
  reg  valid_5; // @[Icache.scala 17:24]
  reg  valid_6; // @[Icache.scala 17:24]
  reg  valid_7; // @[Icache.scala 17:24]
  reg  valid_8; // @[Icache.scala 17:24]
  reg  valid_9; // @[Icache.scala 17:24]
  reg  valid_10; // @[Icache.scala 17:24]
  reg  valid_11; // @[Icache.scala 17:24]
  reg  valid_12; // @[Icache.scala 17:24]
  reg  valid_13; // @[Icache.scala 17:24]
  reg  valid_14; // @[Icache.scala 17:24]
  reg  valid_15; // @[Icache.scala 17:24]
  reg  valid_16; // @[Icache.scala 17:24]
  reg  valid_17; // @[Icache.scala 17:24]
  reg  valid_18; // @[Icache.scala 17:24]
  reg  valid_19; // @[Icache.scala 17:24]
  reg  valid_20; // @[Icache.scala 17:24]
  reg  valid_21; // @[Icache.scala 17:24]
  reg  valid_22; // @[Icache.scala 17:24]
  reg  valid_23; // @[Icache.scala 17:24]
  reg  valid_24; // @[Icache.scala 17:24]
  reg  valid_25; // @[Icache.scala 17:24]
  reg  valid_26; // @[Icache.scala 17:24]
  reg  valid_27; // @[Icache.scala 17:24]
  reg  valid_28; // @[Icache.scala 17:24]
  reg  valid_29; // @[Icache.scala 17:24]
  reg  valid_30; // @[Icache.scala 17:24]
  reg  valid_31; // @[Icache.scala 17:24]
  reg  valid_32; // @[Icache.scala 17:24]
  reg  valid_33; // @[Icache.scala 17:24]
  reg  valid_34; // @[Icache.scala 17:24]
  reg  valid_35; // @[Icache.scala 17:24]
  reg  valid_36; // @[Icache.scala 17:24]
  reg  valid_37; // @[Icache.scala 17:24]
  reg  valid_38; // @[Icache.scala 17:24]
  reg  valid_39; // @[Icache.scala 17:24]
  reg  valid_40; // @[Icache.scala 17:24]
  reg  valid_41; // @[Icache.scala 17:24]
  reg  valid_42; // @[Icache.scala 17:24]
  reg  valid_43; // @[Icache.scala 17:24]
  reg  valid_44; // @[Icache.scala 17:24]
  reg  valid_45; // @[Icache.scala 17:24]
  reg  valid_46; // @[Icache.scala 17:24]
  reg  valid_47; // @[Icache.scala 17:24]
  reg  valid_48; // @[Icache.scala 17:24]
  reg  valid_49; // @[Icache.scala 17:24]
  reg  valid_50; // @[Icache.scala 17:24]
  reg  valid_51; // @[Icache.scala 17:24]
  reg  valid_52; // @[Icache.scala 17:24]
  reg  valid_53; // @[Icache.scala 17:24]
  reg  valid_54; // @[Icache.scala 17:24]
  reg  valid_55; // @[Icache.scala 17:24]
  reg  valid_56; // @[Icache.scala 17:24]
  reg  valid_57; // @[Icache.scala 17:24]
  reg  valid_58; // @[Icache.scala 17:24]
  reg  valid_59; // @[Icache.scala 17:24]
  reg  valid_60; // @[Icache.scala 17:24]
  reg  valid_61; // @[Icache.scala 17:24]
  reg  valid_62; // @[Icache.scala 17:24]
  reg  valid_63; // @[Icache.scala 17:24]
  reg  valid_64; // @[Icache.scala 17:24]
  reg  valid_65; // @[Icache.scala 17:24]
  reg  valid_66; // @[Icache.scala 17:24]
  reg  valid_67; // @[Icache.scala 17:24]
  reg  valid_68; // @[Icache.scala 17:24]
  reg  valid_69; // @[Icache.scala 17:24]
  reg  valid_70; // @[Icache.scala 17:24]
  reg  valid_71; // @[Icache.scala 17:24]
  reg  valid_72; // @[Icache.scala 17:24]
  reg  valid_73; // @[Icache.scala 17:24]
  reg  valid_74; // @[Icache.scala 17:24]
  reg  valid_75; // @[Icache.scala 17:24]
  reg  valid_76; // @[Icache.scala 17:24]
  reg  valid_77; // @[Icache.scala 17:24]
  reg  valid_78; // @[Icache.scala 17:24]
  reg  valid_79; // @[Icache.scala 17:24]
  reg  valid_80; // @[Icache.scala 17:24]
  reg  valid_81; // @[Icache.scala 17:24]
  reg  valid_82; // @[Icache.scala 17:24]
  reg  valid_83; // @[Icache.scala 17:24]
  reg  valid_84; // @[Icache.scala 17:24]
  reg  valid_85; // @[Icache.scala 17:24]
  reg  valid_86; // @[Icache.scala 17:24]
  reg  valid_87; // @[Icache.scala 17:24]
  reg  valid_88; // @[Icache.scala 17:24]
  reg  valid_89; // @[Icache.scala 17:24]
  reg  valid_90; // @[Icache.scala 17:24]
  reg  valid_91; // @[Icache.scala 17:24]
  reg  valid_92; // @[Icache.scala 17:24]
  reg  valid_93; // @[Icache.scala 17:24]
  reg  valid_94; // @[Icache.scala 17:24]
  reg  valid_95; // @[Icache.scala 17:24]
  reg  valid_96; // @[Icache.scala 17:24]
  reg  valid_97; // @[Icache.scala 17:24]
  reg  valid_98; // @[Icache.scala 17:24]
  reg  valid_99; // @[Icache.scala 17:24]
  reg  valid_100; // @[Icache.scala 17:24]
  reg  valid_101; // @[Icache.scala 17:24]
  reg  valid_102; // @[Icache.scala 17:24]
  reg  valid_103; // @[Icache.scala 17:24]
  reg  valid_104; // @[Icache.scala 17:24]
  reg  valid_105; // @[Icache.scala 17:24]
  reg  valid_106; // @[Icache.scala 17:24]
  reg  valid_107; // @[Icache.scala 17:24]
  reg  valid_108; // @[Icache.scala 17:24]
  reg  valid_109; // @[Icache.scala 17:24]
  reg  valid_110; // @[Icache.scala 17:24]
  reg  valid_111; // @[Icache.scala 17:24]
  reg  valid_112; // @[Icache.scala 17:24]
  reg  valid_113; // @[Icache.scala 17:24]
  reg  valid_114; // @[Icache.scala 17:24]
  reg  valid_115; // @[Icache.scala 17:24]
  reg  valid_116; // @[Icache.scala 17:24]
  reg  valid_117; // @[Icache.scala 17:24]
  reg  valid_118; // @[Icache.scala 17:24]
  reg  valid_119; // @[Icache.scala 17:24]
  reg  valid_120; // @[Icache.scala 17:24]
  reg  valid_121; // @[Icache.scala 17:24]
  reg  valid_122; // @[Icache.scala 17:24]
  reg  valid_123; // @[Icache.scala 17:24]
  reg  valid_124; // @[Icache.scala 17:24]
  reg  valid_125; // @[Icache.scala 17:24]
  reg  valid_126; // @[Icache.scala 17:24]
  reg  valid_127; // @[Icache.scala 17:24]
  reg  valid_128; // @[Icache.scala 17:24]
  reg  valid_129; // @[Icache.scala 17:24]
  reg  valid_130; // @[Icache.scala 17:24]
  reg  valid_131; // @[Icache.scala 17:24]
  reg  valid_132; // @[Icache.scala 17:24]
  reg  valid_133; // @[Icache.scala 17:24]
  reg  valid_134; // @[Icache.scala 17:24]
  reg  valid_135; // @[Icache.scala 17:24]
  reg  valid_136; // @[Icache.scala 17:24]
  reg  valid_137; // @[Icache.scala 17:24]
  reg  valid_138; // @[Icache.scala 17:24]
  reg  valid_139; // @[Icache.scala 17:24]
  reg  valid_140; // @[Icache.scala 17:24]
  reg  valid_141; // @[Icache.scala 17:24]
  reg  valid_142; // @[Icache.scala 17:24]
  reg  valid_143; // @[Icache.scala 17:24]
  reg  valid_144; // @[Icache.scala 17:24]
  reg  valid_145; // @[Icache.scala 17:24]
  reg  valid_146; // @[Icache.scala 17:24]
  reg  valid_147; // @[Icache.scala 17:24]
  reg  valid_148; // @[Icache.scala 17:24]
  reg  valid_149; // @[Icache.scala 17:24]
  reg  valid_150; // @[Icache.scala 17:24]
  reg  valid_151; // @[Icache.scala 17:24]
  reg  valid_152; // @[Icache.scala 17:24]
  reg  valid_153; // @[Icache.scala 17:24]
  reg  valid_154; // @[Icache.scala 17:24]
  reg  valid_155; // @[Icache.scala 17:24]
  reg  valid_156; // @[Icache.scala 17:24]
  reg  valid_157; // @[Icache.scala 17:24]
  reg  valid_158; // @[Icache.scala 17:24]
  reg  valid_159; // @[Icache.scala 17:24]
  reg  valid_160; // @[Icache.scala 17:24]
  reg  valid_161; // @[Icache.scala 17:24]
  reg  valid_162; // @[Icache.scala 17:24]
  reg  valid_163; // @[Icache.scala 17:24]
  reg  valid_164; // @[Icache.scala 17:24]
  reg  valid_165; // @[Icache.scala 17:24]
  reg  valid_166; // @[Icache.scala 17:24]
  reg  valid_167; // @[Icache.scala 17:24]
  reg  valid_168; // @[Icache.scala 17:24]
  reg  valid_169; // @[Icache.scala 17:24]
  reg  valid_170; // @[Icache.scala 17:24]
  reg  valid_171; // @[Icache.scala 17:24]
  reg  valid_172; // @[Icache.scala 17:24]
  reg  valid_173; // @[Icache.scala 17:24]
  reg  valid_174; // @[Icache.scala 17:24]
  reg  valid_175; // @[Icache.scala 17:24]
  reg  valid_176; // @[Icache.scala 17:24]
  reg  valid_177; // @[Icache.scala 17:24]
  reg  valid_178; // @[Icache.scala 17:24]
  reg  valid_179; // @[Icache.scala 17:24]
  reg  valid_180; // @[Icache.scala 17:24]
  reg  valid_181; // @[Icache.scala 17:24]
  reg  valid_182; // @[Icache.scala 17:24]
  reg  valid_183; // @[Icache.scala 17:24]
  reg  valid_184; // @[Icache.scala 17:24]
  reg  valid_185; // @[Icache.scala 17:24]
  reg  valid_186; // @[Icache.scala 17:24]
  reg  valid_187; // @[Icache.scala 17:24]
  reg  valid_188; // @[Icache.scala 17:24]
  reg  valid_189; // @[Icache.scala 17:24]
  reg  valid_190; // @[Icache.scala 17:24]
  reg  valid_191; // @[Icache.scala 17:24]
  reg  valid_192; // @[Icache.scala 17:24]
  reg  valid_193; // @[Icache.scala 17:24]
  reg  valid_194; // @[Icache.scala 17:24]
  reg  valid_195; // @[Icache.scala 17:24]
  reg  valid_196; // @[Icache.scala 17:24]
  reg  valid_197; // @[Icache.scala 17:24]
  reg  valid_198; // @[Icache.scala 17:24]
  reg  valid_199; // @[Icache.scala 17:24]
  reg  valid_200; // @[Icache.scala 17:24]
  reg  valid_201; // @[Icache.scala 17:24]
  reg  valid_202; // @[Icache.scala 17:24]
  reg  valid_203; // @[Icache.scala 17:24]
  reg  valid_204; // @[Icache.scala 17:24]
  reg  valid_205; // @[Icache.scala 17:24]
  reg  valid_206; // @[Icache.scala 17:24]
  reg  valid_207; // @[Icache.scala 17:24]
  reg  valid_208; // @[Icache.scala 17:24]
  reg  valid_209; // @[Icache.scala 17:24]
  reg  valid_210; // @[Icache.scala 17:24]
  reg  valid_211; // @[Icache.scala 17:24]
  reg  valid_212; // @[Icache.scala 17:24]
  reg  valid_213; // @[Icache.scala 17:24]
  reg  valid_214; // @[Icache.scala 17:24]
  reg  valid_215; // @[Icache.scala 17:24]
  reg  valid_216; // @[Icache.scala 17:24]
  reg  valid_217; // @[Icache.scala 17:24]
  reg  valid_218; // @[Icache.scala 17:24]
  reg  valid_219; // @[Icache.scala 17:24]
  reg  valid_220; // @[Icache.scala 17:24]
  reg  valid_221; // @[Icache.scala 17:24]
  reg  valid_222; // @[Icache.scala 17:24]
  reg  valid_223; // @[Icache.scala 17:24]
  reg  valid_224; // @[Icache.scala 17:24]
  reg  valid_225; // @[Icache.scala 17:24]
  reg  valid_226; // @[Icache.scala 17:24]
  reg  valid_227; // @[Icache.scala 17:24]
  reg  valid_228; // @[Icache.scala 17:24]
  reg  valid_229; // @[Icache.scala 17:24]
  reg  valid_230; // @[Icache.scala 17:24]
  reg  valid_231; // @[Icache.scala 17:24]
  reg  valid_232; // @[Icache.scala 17:24]
  reg  valid_233; // @[Icache.scala 17:24]
  reg  valid_234; // @[Icache.scala 17:24]
  reg  valid_235; // @[Icache.scala 17:24]
  reg  valid_236; // @[Icache.scala 17:24]
  reg  valid_237; // @[Icache.scala 17:24]
  reg  valid_238; // @[Icache.scala 17:24]
  reg  valid_239; // @[Icache.scala 17:24]
  reg  valid_240; // @[Icache.scala 17:24]
  reg  valid_241; // @[Icache.scala 17:24]
  reg  valid_242; // @[Icache.scala 17:24]
  reg  valid_243; // @[Icache.scala 17:24]
  reg  valid_244; // @[Icache.scala 17:24]
  reg  valid_245; // @[Icache.scala 17:24]
  reg  valid_246; // @[Icache.scala 17:24]
  reg  valid_247; // @[Icache.scala 17:24]
  reg  valid_248; // @[Icache.scala 17:24]
  reg  valid_249; // @[Icache.scala 17:24]
  reg  valid_250; // @[Icache.scala 17:24]
  reg  valid_251; // @[Icache.scala 17:24]
  reg  valid_252; // @[Icache.scala 17:24]
  reg  valid_253; // @[Icache.scala 17:24]
  reg  valid_254; // @[Icache.scala 17:24]
  reg  valid_255; // @[Icache.scala 17:24]
  reg [1:0] state; // @[Icache.scala 25:22]
  reg [31:0] req_addr; // @[Icache.scala 27:27]
  wire  _valid_addr_T = state == 2'h1; // @[Icache.scala 28:30]
  wire [31:0] valid_addr = state == 2'h1 ? io_imem_inst_addr : req_addr; // @[Icache.scala 28:23]
  wire [19:0] req_tag = valid_addr[31:12]; // @[Icache.scala 30:28]
  wire [7:0] req_index = valid_addr[11:4]; // @[Icache.scala 31:28]
  wire [3:0] req_offset = valid_addr[3:0]; // @[Icache.scala 32:28]
  wire [19:0] _GEN_1 = 8'h1 == req_index ? tag_1 : tag_0; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_2 = 8'h2 == req_index ? tag_2 : _GEN_1; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_3 = 8'h3 == req_index ? tag_3 : _GEN_2; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_4 = 8'h4 == req_index ? tag_4 : _GEN_3; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_5 = 8'h5 == req_index ? tag_5 : _GEN_4; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_6 = 8'h6 == req_index ? tag_6 : _GEN_5; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_7 = 8'h7 == req_index ? tag_7 : _GEN_6; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_8 = 8'h8 == req_index ? tag_8 : _GEN_7; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_9 = 8'h9 == req_index ? tag_9 : _GEN_8; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_10 = 8'ha == req_index ? tag_10 : _GEN_9; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_11 = 8'hb == req_index ? tag_11 : _GEN_10; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_12 = 8'hc == req_index ? tag_12 : _GEN_11; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_13 = 8'hd == req_index ? tag_13 : _GEN_12; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_14 = 8'he == req_index ? tag_14 : _GEN_13; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_15 = 8'hf == req_index ? tag_15 : _GEN_14; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_16 = 8'h10 == req_index ? tag_16 : _GEN_15; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_17 = 8'h11 == req_index ? tag_17 : _GEN_16; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_18 = 8'h12 == req_index ? tag_18 : _GEN_17; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_19 = 8'h13 == req_index ? tag_19 : _GEN_18; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_20 = 8'h14 == req_index ? tag_20 : _GEN_19; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_21 = 8'h15 == req_index ? tag_21 : _GEN_20; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_22 = 8'h16 == req_index ? tag_22 : _GEN_21; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_23 = 8'h17 == req_index ? tag_23 : _GEN_22; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_24 = 8'h18 == req_index ? tag_24 : _GEN_23; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_25 = 8'h19 == req_index ? tag_25 : _GEN_24; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_26 = 8'h1a == req_index ? tag_26 : _GEN_25; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_27 = 8'h1b == req_index ? tag_27 : _GEN_26; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_28 = 8'h1c == req_index ? tag_28 : _GEN_27; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_29 = 8'h1d == req_index ? tag_29 : _GEN_28; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_30 = 8'h1e == req_index ? tag_30 : _GEN_29; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_31 = 8'h1f == req_index ? tag_31 : _GEN_30; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_32 = 8'h20 == req_index ? tag_32 : _GEN_31; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_33 = 8'h21 == req_index ? tag_33 : _GEN_32; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_34 = 8'h22 == req_index ? tag_34 : _GEN_33; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_35 = 8'h23 == req_index ? tag_35 : _GEN_34; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_36 = 8'h24 == req_index ? tag_36 : _GEN_35; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_37 = 8'h25 == req_index ? tag_37 : _GEN_36; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_38 = 8'h26 == req_index ? tag_38 : _GEN_37; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_39 = 8'h27 == req_index ? tag_39 : _GEN_38; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_40 = 8'h28 == req_index ? tag_40 : _GEN_39; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_41 = 8'h29 == req_index ? tag_41 : _GEN_40; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_42 = 8'h2a == req_index ? tag_42 : _GEN_41; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_43 = 8'h2b == req_index ? tag_43 : _GEN_42; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_44 = 8'h2c == req_index ? tag_44 : _GEN_43; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_45 = 8'h2d == req_index ? tag_45 : _GEN_44; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_46 = 8'h2e == req_index ? tag_46 : _GEN_45; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_47 = 8'h2f == req_index ? tag_47 : _GEN_46; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_48 = 8'h30 == req_index ? tag_48 : _GEN_47; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_49 = 8'h31 == req_index ? tag_49 : _GEN_48; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_50 = 8'h32 == req_index ? tag_50 : _GEN_49; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_51 = 8'h33 == req_index ? tag_51 : _GEN_50; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_52 = 8'h34 == req_index ? tag_52 : _GEN_51; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_53 = 8'h35 == req_index ? tag_53 : _GEN_52; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_54 = 8'h36 == req_index ? tag_54 : _GEN_53; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_55 = 8'h37 == req_index ? tag_55 : _GEN_54; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_56 = 8'h38 == req_index ? tag_56 : _GEN_55; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_57 = 8'h39 == req_index ? tag_57 : _GEN_56; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_58 = 8'h3a == req_index ? tag_58 : _GEN_57; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_59 = 8'h3b == req_index ? tag_59 : _GEN_58; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_60 = 8'h3c == req_index ? tag_60 : _GEN_59; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_61 = 8'h3d == req_index ? tag_61 : _GEN_60; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_62 = 8'h3e == req_index ? tag_62 : _GEN_61; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_63 = 8'h3f == req_index ? tag_63 : _GEN_62; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_64 = 8'h40 == req_index ? tag_64 : _GEN_63; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_65 = 8'h41 == req_index ? tag_65 : _GEN_64; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_66 = 8'h42 == req_index ? tag_66 : _GEN_65; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_67 = 8'h43 == req_index ? tag_67 : _GEN_66; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_68 = 8'h44 == req_index ? tag_68 : _GEN_67; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_69 = 8'h45 == req_index ? tag_69 : _GEN_68; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_70 = 8'h46 == req_index ? tag_70 : _GEN_69; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_71 = 8'h47 == req_index ? tag_71 : _GEN_70; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_72 = 8'h48 == req_index ? tag_72 : _GEN_71; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_73 = 8'h49 == req_index ? tag_73 : _GEN_72; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_74 = 8'h4a == req_index ? tag_74 : _GEN_73; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_75 = 8'h4b == req_index ? tag_75 : _GEN_74; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_76 = 8'h4c == req_index ? tag_76 : _GEN_75; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_77 = 8'h4d == req_index ? tag_77 : _GEN_76; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_78 = 8'h4e == req_index ? tag_78 : _GEN_77; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_79 = 8'h4f == req_index ? tag_79 : _GEN_78; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_80 = 8'h50 == req_index ? tag_80 : _GEN_79; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_81 = 8'h51 == req_index ? tag_81 : _GEN_80; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_82 = 8'h52 == req_index ? tag_82 : _GEN_81; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_83 = 8'h53 == req_index ? tag_83 : _GEN_82; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_84 = 8'h54 == req_index ? tag_84 : _GEN_83; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_85 = 8'h55 == req_index ? tag_85 : _GEN_84; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_86 = 8'h56 == req_index ? tag_86 : _GEN_85; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_87 = 8'h57 == req_index ? tag_87 : _GEN_86; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_88 = 8'h58 == req_index ? tag_88 : _GEN_87; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_89 = 8'h59 == req_index ? tag_89 : _GEN_88; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_90 = 8'h5a == req_index ? tag_90 : _GEN_89; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_91 = 8'h5b == req_index ? tag_91 : _GEN_90; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_92 = 8'h5c == req_index ? tag_92 : _GEN_91; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_93 = 8'h5d == req_index ? tag_93 : _GEN_92; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_94 = 8'h5e == req_index ? tag_94 : _GEN_93; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_95 = 8'h5f == req_index ? tag_95 : _GEN_94; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_96 = 8'h60 == req_index ? tag_96 : _GEN_95; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_97 = 8'h61 == req_index ? tag_97 : _GEN_96; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_98 = 8'h62 == req_index ? tag_98 : _GEN_97; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_99 = 8'h63 == req_index ? tag_99 : _GEN_98; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_100 = 8'h64 == req_index ? tag_100 : _GEN_99; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_101 = 8'h65 == req_index ? tag_101 : _GEN_100; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_102 = 8'h66 == req_index ? tag_102 : _GEN_101; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_103 = 8'h67 == req_index ? tag_103 : _GEN_102; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_104 = 8'h68 == req_index ? tag_104 : _GEN_103; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_105 = 8'h69 == req_index ? tag_105 : _GEN_104; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_106 = 8'h6a == req_index ? tag_106 : _GEN_105; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_107 = 8'h6b == req_index ? tag_107 : _GEN_106; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_108 = 8'h6c == req_index ? tag_108 : _GEN_107; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_109 = 8'h6d == req_index ? tag_109 : _GEN_108; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_110 = 8'h6e == req_index ? tag_110 : _GEN_109; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_111 = 8'h6f == req_index ? tag_111 : _GEN_110; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_112 = 8'h70 == req_index ? tag_112 : _GEN_111; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_113 = 8'h71 == req_index ? tag_113 : _GEN_112; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_114 = 8'h72 == req_index ? tag_114 : _GEN_113; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_115 = 8'h73 == req_index ? tag_115 : _GEN_114; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_116 = 8'h74 == req_index ? tag_116 : _GEN_115; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_117 = 8'h75 == req_index ? tag_117 : _GEN_116; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_118 = 8'h76 == req_index ? tag_118 : _GEN_117; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_119 = 8'h77 == req_index ? tag_119 : _GEN_118; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_120 = 8'h78 == req_index ? tag_120 : _GEN_119; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_121 = 8'h79 == req_index ? tag_121 : _GEN_120; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_122 = 8'h7a == req_index ? tag_122 : _GEN_121; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_123 = 8'h7b == req_index ? tag_123 : _GEN_122; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_124 = 8'h7c == req_index ? tag_124 : _GEN_123; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_125 = 8'h7d == req_index ? tag_125 : _GEN_124; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_126 = 8'h7e == req_index ? tag_126 : _GEN_125; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_127 = 8'h7f == req_index ? tag_127 : _GEN_126; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_128 = 8'h80 == req_index ? tag_128 : _GEN_127; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_129 = 8'h81 == req_index ? tag_129 : _GEN_128; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_130 = 8'h82 == req_index ? tag_130 : _GEN_129; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_131 = 8'h83 == req_index ? tag_131 : _GEN_130; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_132 = 8'h84 == req_index ? tag_132 : _GEN_131; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_133 = 8'h85 == req_index ? tag_133 : _GEN_132; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_134 = 8'h86 == req_index ? tag_134 : _GEN_133; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_135 = 8'h87 == req_index ? tag_135 : _GEN_134; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_136 = 8'h88 == req_index ? tag_136 : _GEN_135; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_137 = 8'h89 == req_index ? tag_137 : _GEN_136; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_138 = 8'h8a == req_index ? tag_138 : _GEN_137; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_139 = 8'h8b == req_index ? tag_139 : _GEN_138; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_140 = 8'h8c == req_index ? tag_140 : _GEN_139; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_141 = 8'h8d == req_index ? tag_141 : _GEN_140; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_142 = 8'h8e == req_index ? tag_142 : _GEN_141; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_143 = 8'h8f == req_index ? tag_143 : _GEN_142; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_144 = 8'h90 == req_index ? tag_144 : _GEN_143; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_145 = 8'h91 == req_index ? tag_145 : _GEN_144; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_146 = 8'h92 == req_index ? tag_146 : _GEN_145; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_147 = 8'h93 == req_index ? tag_147 : _GEN_146; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_148 = 8'h94 == req_index ? tag_148 : _GEN_147; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_149 = 8'h95 == req_index ? tag_149 : _GEN_148; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_150 = 8'h96 == req_index ? tag_150 : _GEN_149; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_151 = 8'h97 == req_index ? tag_151 : _GEN_150; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_152 = 8'h98 == req_index ? tag_152 : _GEN_151; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_153 = 8'h99 == req_index ? tag_153 : _GEN_152; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_154 = 8'h9a == req_index ? tag_154 : _GEN_153; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_155 = 8'h9b == req_index ? tag_155 : _GEN_154; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_156 = 8'h9c == req_index ? tag_156 : _GEN_155; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_157 = 8'h9d == req_index ? tag_157 : _GEN_156; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_158 = 8'h9e == req_index ? tag_158 : _GEN_157; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_159 = 8'h9f == req_index ? tag_159 : _GEN_158; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_160 = 8'ha0 == req_index ? tag_160 : _GEN_159; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_161 = 8'ha1 == req_index ? tag_161 : _GEN_160; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_162 = 8'ha2 == req_index ? tag_162 : _GEN_161; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_163 = 8'ha3 == req_index ? tag_163 : _GEN_162; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_164 = 8'ha4 == req_index ? tag_164 : _GEN_163; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_165 = 8'ha5 == req_index ? tag_165 : _GEN_164; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_166 = 8'ha6 == req_index ? tag_166 : _GEN_165; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_167 = 8'ha7 == req_index ? tag_167 : _GEN_166; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_168 = 8'ha8 == req_index ? tag_168 : _GEN_167; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_169 = 8'ha9 == req_index ? tag_169 : _GEN_168; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_170 = 8'haa == req_index ? tag_170 : _GEN_169; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_171 = 8'hab == req_index ? tag_171 : _GEN_170; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_172 = 8'hac == req_index ? tag_172 : _GEN_171; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_173 = 8'had == req_index ? tag_173 : _GEN_172; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_174 = 8'hae == req_index ? tag_174 : _GEN_173; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_175 = 8'haf == req_index ? tag_175 : _GEN_174; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_176 = 8'hb0 == req_index ? tag_176 : _GEN_175; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_177 = 8'hb1 == req_index ? tag_177 : _GEN_176; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_178 = 8'hb2 == req_index ? tag_178 : _GEN_177; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_179 = 8'hb3 == req_index ? tag_179 : _GEN_178; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_180 = 8'hb4 == req_index ? tag_180 : _GEN_179; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_181 = 8'hb5 == req_index ? tag_181 : _GEN_180; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_182 = 8'hb6 == req_index ? tag_182 : _GEN_181; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_183 = 8'hb7 == req_index ? tag_183 : _GEN_182; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_184 = 8'hb8 == req_index ? tag_184 : _GEN_183; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_185 = 8'hb9 == req_index ? tag_185 : _GEN_184; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_186 = 8'hba == req_index ? tag_186 : _GEN_185; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_187 = 8'hbb == req_index ? tag_187 : _GEN_186; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_188 = 8'hbc == req_index ? tag_188 : _GEN_187; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_189 = 8'hbd == req_index ? tag_189 : _GEN_188; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_190 = 8'hbe == req_index ? tag_190 : _GEN_189; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_191 = 8'hbf == req_index ? tag_191 : _GEN_190; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_192 = 8'hc0 == req_index ? tag_192 : _GEN_191; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_193 = 8'hc1 == req_index ? tag_193 : _GEN_192; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_194 = 8'hc2 == req_index ? tag_194 : _GEN_193; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_195 = 8'hc3 == req_index ? tag_195 : _GEN_194; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_196 = 8'hc4 == req_index ? tag_196 : _GEN_195; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_197 = 8'hc5 == req_index ? tag_197 : _GEN_196; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_198 = 8'hc6 == req_index ? tag_198 : _GEN_197; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_199 = 8'hc7 == req_index ? tag_199 : _GEN_198; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_200 = 8'hc8 == req_index ? tag_200 : _GEN_199; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_201 = 8'hc9 == req_index ? tag_201 : _GEN_200; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_202 = 8'hca == req_index ? tag_202 : _GEN_201; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_203 = 8'hcb == req_index ? tag_203 : _GEN_202; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_204 = 8'hcc == req_index ? tag_204 : _GEN_203; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_205 = 8'hcd == req_index ? tag_205 : _GEN_204; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_206 = 8'hce == req_index ? tag_206 : _GEN_205; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_207 = 8'hcf == req_index ? tag_207 : _GEN_206; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_208 = 8'hd0 == req_index ? tag_208 : _GEN_207; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_209 = 8'hd1 == req_index ? tag_209 : _GEN_208; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_210 = 8'hd2 == req_index ? tag_210 : _GEN_209; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_211 = 8'hd3 == req_index ? tag_211 : _GEN_210; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_212 = 8'hd4 == req_index ? tag_212 : _GEN_211; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_213 = 8'hd5 == req_index ? tag_213 : _GEN_212; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_214 = 8'hd6 == req_index ? tag_214 : _GEN_213; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_215 = 8'hd7 == req_index ? tag_215 : _GEN_214; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_216 = 8'hd8 == req_index ? tag_216 : _GEN_215; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_217 = 8'hd9 == req_index ? tag_217 : _GEN_216; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_218 = 8'hda == req_index ? tag_218 : _GEN_217; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_219 = 8'hdb == req_index ? tag_219 : _GEN_218; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_220 = 8'hdc == req_index ? tag_220 : _GEN_219; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_221 = 8'hdd == req_index ? tag_221 : _GEN_220; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_222 = 8'hde == req_index ? tag_222 : _GEN_221; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_223 = 8'hdf == req_index ? tag_223 : _GEN_222; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_224 = 8'he0 == req_index ? tag_224 : _GEN_223; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_225 = 8'he1 == req_index ? tag_225 : _GEN_224; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_226 = 8'he2 == req_index ? tag_226 : _GEN_225; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_227 = 8'he3 == req_index ? tag_227 : _GEN_226; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_228 = 8'he4 == req_index ? tag_228 : _GEN_227; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_229 = 8'he5 == req_index ? tag_229 : _GEN_228; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_230 = 8'he6 == req_index ? tag_230 : _GEN_229; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_231 = 8'he7 == req_index ? tag_231 : _GEN_230; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_232 = 8'he8 == req_index ? tag_232 : _GEN_231; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_233 = 8'he9 == req_index ? tag_233 : _GEN_232; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_234 = 8'hea == req_index ? tag_234 : _GEN_233; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_235 = 8'heb == req_index ? tag_235 : _GEN_234; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_236 = 8'hec == req_index ? tag_236 : _GEN_235; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_237 = 8'hed == req_index ? tag_237 : _GEN_236; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_238 = 8'hee == req_index ? tag_238 : _GEN_237; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_239 = 8'hef == req_index ? tag_239 : _GEN_238; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_240 = 8'hf0 == req_index ? tag_240 : _GEN_239; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_241 = 8'hf1 == req_index ? tag_241 : _GEN_240; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_242 = 8'hf2 == req_index ? tag_242 : _GEN_241; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_243 = 8'hf3 == req_index ? tag_243 : _GEN_242; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_244 = 8'hf4 == req_index ? tag_244 : _GEN_243; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_245 = 8'hf5 == req_index ? tag_245 : _GEN_244; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_246 = 8'hf6 == req_index ? tag_246 : _GEN_245; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_247 = 8'hf7 == req_index ? tag_247 : _GEN_246; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_248 = 8'hf8 == req_index ? tag_248 : _GEN_247; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_249 = 8'hf9 == req_index ? tag_249 : _GEN_248; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_250 = 8'hfa == req_index ? tag_250 : _GEN_249; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_251 = 8'hfb == req_index ? tag_251 : _GEN_250; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_252 = 8'hfc == req_index ? tag_252 : _GEN_251; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_253 = 8'hfd == req_index ? tag_253 : _GEN_252; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_254 = 8'hfe == req_index ? tag_254 : _GEN_253; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire [19:0] _GEN_255 = 8'hff == req_index ? tag_255 : _GEN_254; // @[Icache.scala 35:32 Icache.scala 35:32]
  wire  _GEN_257 = 8'h1 == req_index ? valid_1 : valid_0; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_258 = 8'h2 == req_index ? valid_2 : _GEN_257; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_259 = 8'h3 == req_index ? valid_3 : _GEN_258; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_260 = 8'h4 == req_index ? valid_4 : _GEN_259; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_261 = 8'h5 == req_index ? valid_5 : _GEN_260; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_262 = 8'h6 == req_index ? valid_6 : _GEN_261; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_263 = 8'h7 == req_index ? valid_7 : _GEN_262; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_264 = 8'h8 == req_index ? valid_8 : _GEN_263; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_265 = 8'h9 == req_index ? valid_9 : _GEN_264; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_266 = 8'ha == req_index ? valid_10 : _GEN_265; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_267 = 8'hb == req_index ? valid_11 : _GEN_266; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_268 = 8'hc == req_index ? valid_12 : _GEN_267; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_269 = 8'hd == req_index ? valid_13 : _GEN_268; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_270 = 8'he == req_index ? valid_14 : _GEN_269; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_271 = 8'hf == req_index ? valid_15 : _GEN_270; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_272 = 8'h10 == req_index ? valid_16 : _GEN_271; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_273 = 8'h11 == req_index ? valid_17 : _GEN_272; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_274 = 8'h12 == req_index ? valid_18 : _GEN_273; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_275 = 8'h13 == req_index ? valid_19 : _GEN_274; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_276 = 8'h14 == req_index ? valid_20 : _GEN_275; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_277 = 8'h15 == req_index ? valid_21 : _GEN_276; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_278 = 8'h16 == req_index ? valid_22 : _GEN_277; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_279 = 8'h17 == req_index ? valid_23 : _GEN_278; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_280 = 8'h18 == req_index ? valid_24 : _GEN_279; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_281 = 8'h19 == req_index ? valid_25 : _GEN_280; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_282 = 8'h1a == req_index ? valid_26 : _GEN_281; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_283 = 8'h1b == req_index ? valid_27 : _GEN_282; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_284 = 8'h1c == req_index ? valid_28 : _GEN_283; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_285 = 8'h1d == req_index ? valid_29 : _GEN_284; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_286 = 8'h1e == req_index ? valid_30 : _GEN_285; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_287 = 8'h1f == req_index ? valid_31 : _GEN_286; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_288 = 8'h20 == req_index ? valid_32 : _GEN_287; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_289 = 8'h21 == req_index ? valid_33 : _GEN_288; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_290 = 8'h22 == req_index ? valid_34 : _GEN_289; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_291 = 8'h23 == req_index ? valid_35 : _GEN_290; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_292 = 8'h24 == req_index ? valid_36 : _GEN_291; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_293 = 8'h25 == req_index ? valid_37 : _GEN_292; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_294 = 8'h26 == req_index ? valid_38 : _GEN_293; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_295 = 8'h27 == req_index ? valid_39 : _GEN_294; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_296 = 8'h28 == req_index ? valid_40 : _GEN_295; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_297 = 8'h29 == req_index ? valid_41 : _GEN_296; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_298 = 8'h2a == req_index ? valid_42 : _GEN_297; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_299 = 8'h2b == req_index ? valid_43 : _GEN_298; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_300 = 8'h2c == req_index ? valid_44 : _GEN_299; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_301 = 8'h2d == req_index ? valid_45 : _GEN_300; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_302 = 8'h2e == req_index ? valid_46 : _GEN_301; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_303 = 8'h2f == req_index ? valid_47 : _GEN_302; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_304 = 8'h30 == req_index ? valid_48 : _GEN_303; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_305 = 8'h31 == req_index ? valid_49 : _GEN_304; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_306 = 8'h32 == req_index ? valid_50 : _GEN_305; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_307 = 8'h33 == req_index ? valid_51 : _GEN_306; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_308 = 8'h34 == req_index ? valid_52 : _GEN_307; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_309 = 8'h35 == req_index ? valid_53 : _GEN_308; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_310 = 8'h36 == req_index ? valid_54 : _GEN_309; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_311 = 8'h37 == req_index ? valid_55 : _GEN_310; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_312 = 8'h38 == req_index ? valid_56 : _GEN_311; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_313 = 8'h39 == req_index ? valid_57 : _GEN_312; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_314 = 8'h3a == req_index ? valid_58 : _GEN_313; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_315 = 8'h3b == req_index ? valid_59 : _GEN_314; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_316 = 8'h3c == req_index ? valid_60 : _GEN_315; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_317 = 8'h3d == req_index ? valid_61 : _GEN_316; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_318 = 8'h3e == req_index ? valid_62 : _GEN_317; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_319 = 8'h3f == req_index ? valid_63 : _GEN_318; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_320 = 8'h40 == req_index ? valid_64 : _GEN_319; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_321 = 8'h41 == req_index ? valid_65 : _GEN_320; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_322 = 8'h42 == req_index ? valid_66 : _GEN_321; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_323 = 8'h43 == req_index ? valid_67 : _GEN_322; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_324 = 8'h44 == req_index ? valid_68 : _GEN_323; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_325 = 8'h45 == req_index ? valid_69 : _GEN_324; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_326 = 8'h46 == req_index ? valid_70 : _GEN_325; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_327 = 8'h47 == req_index ? valid_71 : _GEN_326; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_328 = 8'h48 == req_index ? valid_72 : _GEN_327; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_329 = 8'h49 == req_index ? valid_73 : _GEN_328; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_330 = 8'h4a == req_index ? valid_74 : _GEN_329; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_331 = 8'h4b == req_index ? valid_75 : _GEN_330; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_332 = 8'h4c == req_index ? valid_76 : _GEN_331; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_333 = 8'h4d == req_index ? valid_77 : _GEN_332; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_334 = 8'h4e == req_index ? valid_78 : _GEN_333; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_335 = 8'h4f == req_index ? valid_79 : _GEN_334; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_336 = 8'h50 == req_index ? valid_80 : _GEN_335; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_337 = 8'h51 == req_index ? valid_81 : _GEN_336; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_338 = 8'h52 == req_index ? valid_82 : _GEN_337; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_339 = 8'h53 == req_index ? valid_83 : _GEN_338; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_340 = 8'h54 == req_index ? valid_84 : _GEN_339; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_341 = 8'h55 == req_index ? valid_85 : _GEN_340; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_342 = 8'h56 == req_index ? valid_86 : _GEN_341; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_343 = 8'h57 == req_index ? valid_87 : _GEN_342; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_344 = 8'h58 == req_index ? valid_88 : _GEN_343; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_345 = 8'h59 == req_index ? valid_89 : _GEN_344; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_346 = 8'h5a == req_index ? valid_90 : _GEN_345; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_347 = 8'h5b == req_index ? valid_91 : _GEN_346; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_348 = 8'h5c == req_index ? valid_92 : _GEN_347; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_349 = 8'h5d == req_index ? valid_93 : _GEN_348; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_350 = 8'h5e == req_index ? valid_94 : _GEN_349; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_351 = 8'h5f == req_index ? valid_95 : _GEN_350; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_352 = 8'h60 == req_index ? valid_96 : _GEN_351; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_353 = 8'h61 == req_index ? valid_97 : _GEN_352; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_354 = 8'h62 == req_index ? valid_98 : _GEN_353; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_355 = 8'h63 == req_index ? valid_99 : _GEN_354; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_356 = 8'h64 == req_index ? valid_100 : _GEN_355; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_357 = 8'h65 == req_index ? valid_101 : _GEN_356; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_358 = 8'h66 == req_index ? valid_102 : _GEN_357; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_359 = 8'h67 == req_index ? valid_103 : _GEN_358; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_360 = 8'h68 == req_index ? valid_104 : _GEN_359; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_361 = 8'h69 == req_index ? valid_105 : _GEN_360; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_362 = 8'h6a == req_index ? valid_106 : _GEN_361; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_363 = 8'h6b == req_index ? valid_107 : _GEN_362; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_364 = 8'h6c == req_index ? valid_108 : _GEN_363; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_365 = 8'h6d == req_index ? valid_109 : _GEN_364; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_366 = 8'h6e == req_index ? valid_110 : _GEN_365; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_367 = 8'h6f == req_index ? valid_111 : _GEN_366; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_368 = 8'h70 == req_index ? valid_112 : _GEN_367; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_369 = 8'h71 == req_index ? valid_113 : _GEN_368; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_370 = 8'h72 == req_index ? valid_114 : _GEN_369; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_371 = 8'h73 == req_index ? valid_115 : _GEN_370; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_372 = 8'h74 == req_index ? valid_116 : _GEN_371; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_373 = 8'h75 == req_index ? valid_117 : _GEN_372; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_374 = 8'h76 == req_index ? valid_118 : _GEN_373; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_375 = 8'h77 == req_index ? valid_119 : _GEN_374; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_376 = 8'h78 == req_index ? valid_120 : _GEN_375; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_377 = 8'h79 == req_index ? valid_121 : _GEN_376; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_378 = 8'h7a == req_index ? valid_122 : _GEN_377; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_379 = 8'h7b == req_index ? valid_123 : _GEN_378; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_380 = 8'h7c == req_index ? valid_124 : _GEN_379; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_381 = 8'h7d == req_index ? valid_125 : _GEN_380; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_382 = 8'h7e == req_index ? valid_126 : _GEN_381; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_383 = 8'h7f == req_index ? valid_127 : _GEN_382; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_384 = 8'h80 == req_index ? valid_128 : _GEN_383; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_385 = 8'h81 == req_index ? valid_129 : _GEN_384; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_386 = 8'h82 == req_index ? valid_130 : _GEN_385; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_387 = 8'h83 == req_index ? valid_131 : _GEN_386; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_388 = 8'h84 == req_index ? valid_132 : _GEN_387; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_389 = 8'h85 == req_index ? valid_133 : _GEN_388; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_390 = 8'h86 == req_index ? valid_134 : _GEN_389; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_391 = 8'h87 == req_index ? valid_135 : _GEN_390; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_392 = 8'h88 == req_index ? valid_136 : _GEN_391; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_393 = 8'h89 == req_index ? valid_137 : _GEN_392; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_394 = 8'h8a == req_index ? valid_138 : _GEN_393; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_395 = 8'h8b == req_index ? valid_139 : _GEN_394; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_396 = 8'h8c == req_index ? valid_140 : _GEN_395; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_397 = 8'h8d == req_index ? valid_141 : _GEN_396; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_398 = 8'h8e == req_index ? valid_142 : _GEN_397; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_399 = 8'h8f == req_index ? valid_143 : _GEN_398; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_400 = 8'h90 == req_index ? valid_144 : _GEN_399; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_401 = 8'h91 == req_index ? valid_145 : _GEN_400; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_402 = 8'h92 == req_index ? valid_146 : _GEN_401; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_403 = 8'h93 == req_index ? valid_147 : _GEN_402; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_404 = 8'h94 == req_index ? valid_148 : _GEN_403; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_405 = 8'h95 == req_index ? valid_149 : _GEN_404; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_406 = 8'h96 == req_index ? valid_150 : _GEN_405; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_407 = 8'h97 == req_index ? valid_151 : _GEN_406; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_408 = 8'h98 == req_index ? valid_152 : _GEN_407; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_409 = 8'h99 == req_index ? valid_153 : _GEN_408; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_410 = 8'h9a == req_index ? valid_154 : _GEN_409; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_411 = 8'h9b == req_index ? valid_155 : _GEN_410; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_412 = 8'h9c == req_index ? valid_156 : _GEN_411; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_413 = 8'h9d == req_index ? valid_157 : _GEN_412; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_414 = 8'h9e == req_index ? valid_158 : _GEN_413; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_415 = 8'h9f == req_index ? valid_159 : _GEN_414; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_416 = 8'ha0 == req_index ? valid_160 : _GEN_415; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_417 = 8'ha1 == req_index ? valid_161 : _GEN_416; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_418 = 8'ha2 == req_index ? valid_162 : _GEN_417; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_419 = 8'ha3 == req_index ? valid_163 : _GEN_418; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_420 = 8'ha4 == req_index ? valid_164 : _GEN_419; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_421 = 8'ha5 == req_index ? valid_165 : _GEN_420; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_422 = 8'ha6 == req_index ? valid_166 : _GEN_421; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_423 = 8'ha7 == req_index ? valid_167 : _GEN_422; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_424 = 8'ha8 == req_index ? valid_168 : _GEN_423; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_425 = 8'ha9 == req_index ? valid_169 : _GEN_424; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_426 = 8'haa == req_index ? valid_170 : _GEN_425; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_427 = 8'hab == req_index ? valid_171 : _GEN_426; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_428 = 8'hac == req_index ? valid_172 : _GEN_427; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_429 = 8'had == req_index ? valid_173 : _GEN_428; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_430 = 8'hae == req_index ? valid_174 : _GEN_429; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_431 = 8'haf == req_index ? valid_175 : _GEN_430; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_432 = 8'hb0 == req_index ? valid_176 : _GEN_431; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_433 = 8'hb1 == req_index ? valid_177 : _GEN_432; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_434 = 8'hb2 == req_index ? valid_178 : _GEN_433; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_435 = 8'hb3 == req_index ? valid_179 : _GEN_434; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_436 = 8'hb4 == req_index ? valid_180 : _GEN_435; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_437 = 8'hb5 == req_index ? valid_181 : _GEN_436; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_438 = 8'hb6 == req_index ? valid_182 : _GEN_437; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_439 = 8'hb7 == req_index ? valid_183 : _GEN_438; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_440 = 8'hb8 == req_index ? valid_184 : _GEN_439; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_441 = 8'hb9 == req_index ? valid_185 : _GEN_440; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_442 = 8'hba == req_index ? valid_186 : _GEN_441; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_443 = 8'hbb == req_index ? valid_187 : _GEN_442; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_444 = 8'hbc == req_index ? valid_188 : _GEN_443; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_445 = 8'hbd == req_index ? valid_189 : _GEN_444; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_446 = 8'hbe == req_index ? valid_190 : _GEN_445; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_447 = 8'hbf == req_index ? valid_191 : _GEN_446; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_448 = 8'hc0 == req_index ? valid_192 : _GEN_447; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_449 = 8'hc1 == req_index ? valid_193 : _GEN_448; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_450 = 8'hc2 == req_index ? valid_194 : _GEN_449; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_451 = 8'hc3 == req_index ? valid_195 : _GEN_450; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_452 = 8'hc4 == req_index ? valid_196 : _GEN_451; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_453 = 8'hc5 == req_index ? valid_197 : _GEN_452; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_454 = 8'hc6 == req_index ? valid_198 : _GEN_453; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_455 = 8'hc7 == req_index ? valid_199 : _GEN_454; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_456 = 8'hc8 == req_index ? valid_200 : _GEN_455; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_457 = 8'hc9 == req_index ? valid_201 : _GEN_456; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_458 = 8'hca == req_index ? valid_202 : _GEN_457; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_459 = 8'hcb == req_index ? valid_203 : _GEN_458; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_460 = 8'hcc == req_index ? valid_204 : _GEN_459; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_461 = 8'hcd == req_index ? valid_205 : _GEN_460; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_462 = 8'hce == req_index ? valid_206 : _GEN_461; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_463 = 8'hcf == req_index ? valid_207 : _GEN_462; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_464 = 8'hd0 == req_index ? valid_208 : _GEN_463; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_465 = 8'hd1 == req_index ? valid_209 : _GEN_464; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_466 = 8'hd2 == req_index ? valid_210 : _GEN_465; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_467 = 8'hd3 == req_index ? valid_211 : _GEN_466; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_468 = 8'hd4 == req_index ? valid_212 : _GEN_467; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_469 = 8'hd5 == req_index ? valid_213 : _GEN_468; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_470 = 8'hd6 == req_index ? valid_214 : _GEN_469; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_471 = 8'hd7 == req_index ? valid_215 : _GEN_470; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_472 = 8'hd8 == req_index ? valid_216 : _GEN_471; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_473 = 8'hd9 == req_index ? valid_217 : _GEN_472; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_474 = 8'hda == req_index ? valid_218 : _GEN_473; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_475 = 8'hdb == req_index ? valid_219 : _GEN_474; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_476 = 8'hdc == req_index ? valid_220 : _GEN_475; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_477 = 8'hdd == req_index ? valid_221 : _GEN_476; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_478 = 8'hde == req_index ? valid_222 : _GEN_477; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_479 = 8'hdf == req_index ? valid_223 : _GEN_478; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_480 = 8'he0 == req_index ? valid_224 : _GEN_479; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_481 = 8'he1 == req_index ? valid_225 : _GEN_480; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_482 = 8'he2 == req_index ? valid_226 : _GEN_481; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_483 = 8'he3 == req_index ? valid_227 : _GEN_482; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_484 = 8'he4 == req_index ? valid_228 : _GEN_483; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_485 = 8'he5 == req_index ? valid_229 : _GEN_484; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_486 = 8'he6 == req_index ? valid_230 : _GEN_485; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_487 = 8'he7 == req_index ? valid_231 : _GEN_486; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_488 = 8'he8 == req_index ? valid_232 : _GEN_487; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_489 = 8'he9 == req_index ? valid_233 : _GEN_488; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_490 = 8'hea == req_index ? valid_234 : _GEN_489; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_491 = 8'heb == req_index ? valid_235 : _GEN_490; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_492 = 8'hec == req_index ? valid_236 : _GEN_491; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_493 = 8'hed == req_index ? valid_237 : _GEN_492; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_494 = 8'hee == req_index ? valid_238 : _GEN_493; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_495 = 8'hef == req_index ? valid_239 : _GEN_494; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_496 = 8'hf0 == req_index ? valid_240 : _GEN_495; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_497 = 8'hf1 == req_index ? valid_241 : _GEN_496; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_498 = 8'hf2 == req_index ? valid_242 : _GEN_497; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_499 = 8'hf3 == req_index ? valid_243 : _GEN_498; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_500 = 8'hf4 == req_index ? valid_244 : _GEN_499; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_501 = 8'hf5 == req_index ? valid_245 : _GEN_500; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_502 = 8'hf6 == req_index ? valid_246 : _GEN_501; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_503 = 8'hf7 == req_index ? valid_247 : _GEN_502; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_504 = 8'hf8 == req_index ? valid_248 : _GEN_503; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_505 = 8'hf9 == req_index ? valid_249 : _GEN_504; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_506 = 8'hfa == req_index ? valid_250 : _GEN_505; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_507 = 8'hfb == req_index ? valid_251 : _GEN_506; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_508 = 8'hfc == req_index ? valid_252 : _GEN_507; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_509 = 8'hfd == req_index ? valid_253 : _GEN_508; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_510 = 8'hfe == req_index ? valid_254 : _GEN_509; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  _GEN_511 = 8'hff == req_index ? valid_255 : _GEN_510; // @[Icache.scala 35:45 Icache.scala 35:45]
  wire  cache_hit = _GEN_255 == req_tag & _GEN_511; // @[Icache.scala 35:45]
  wire [127:0] cache_data_out = req_Q; // @[Icache.scala 37:28 Icache.scala 120:18]
  wire [31:0] _inst_read_T_6 = 2'h1 == req_offset[3:2] ? cache_data_out[63:32] : cache_data_out[31:0]; // @[Mux.scala 80:57]
  wire [31:0] _inst_read_T_8 = 2'h2 == req_offset[3:2] ? cache_data_out[95:64] : _inst_read_T_6; // @[Mux.scala 80:57]
  reg  cache_fill; // @[Icache.scala 51:28]
  reg  cache_wen; // @[Icache.scala 52:28]
  reg [127:0] cache_wdata; // @[Icache.scala 53:28]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_514 = cache_hit ? 2'h1 : 2'h2; // @[Icache.scala 64:26 Icache.scala 66:20 Icache.scala 70:20]
  wire  _T_2 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = ~cache_fill; // @[Icache.scala 79:13]
  wire [1:0] _GEN_517 = ~cache_fill ? 2'h2 : 2'h3; // @[Icache.scala 79:26 Icache.scala 80:21 Icache.scala 87:21]
  wire [31:0] _GEN_520 = ~cache_fill ? req_addr : 32'h0; // @[Icache.scala 79:26 Icache.scala 83:21]
  wire  _GEN_522 = io_out_inst_ready | cache_fill; // @[Icache.scala 89:29 Icache.scala 90:21 Icache.scala 51:28]
  wire  _GEN_523 = io_out_inst_ready | cache_wen; // @[Icache.scala 89:29 Icache.scala 91:21 Icache.scala 52:28]
  wire [127:0] _GEN_524 = io_out_inst_ready ? io_out_inst_read : cache_wdata; // @[Icache.scala 89:29 Icache.scala 92:21 Icache.scala 53:28]
  wire  _GEN_525 = io_out_inst_ready ? 1'h0 : _T_3; // @[Icache.scala 89:29 Icache.scala 93:21]
  wire  _T_4 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire  _GEN_526 = 8'h0 == req_index | valid_0; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_527 = 8'h1 == req_index | valid_1; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_528 = 8'h2 == req_index | valid_2; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_529 = 8'h3 == req_index | valid_3; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_530 = 8'h4 == req_index | valid_4; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_531 = 8'h5 == req_index | valid_5; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_532 = 8'h6 == req_index | valid_6; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_533 = 8'h7 == req_index | valid_7; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_534 = 8'h8 == req_index | valid_8; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_535 = 8'h9 == req_index | valid_9; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_536 = 8'ha == req_index | valid_10; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_537 = 8'hb == req_index | valid_11; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_538 = 8'hc == req_index | valid_12; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_539 = 8'hd == req_index | valid_13; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_540 = 8'he == req_index | valid_14; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_541 = 8'hf == req_index | valid_15; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_542 = 8'h10 == req_index | valid_16; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_543 = 8'h11 == req_index | valid_17; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_544 = 8'h12 == req_index | valid_18; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_545 = 8'h13 == req_index | valid_19; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_546 = 8'h14 == req_index | valid_20; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_547 = 8'h15 == req_index | valid_21; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_548 = 8'h16 == req_index | valid_22; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_549 = 8'h17 == req_index | valid_23; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_550 = 8'h18 == req_index | valid_24; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_551 = 8'h19 == req_index | valid_25; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_552 = 8'h1a == req_index | valid_26; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_553 = 8'h1b == req_index | valid_27; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_554 = 8'h1c == req_index | valid_28; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_555 = 8'h1d == req_index | valid_29; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_556 = 8'h1e == req_index | valid_30; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_557 = 8'h1f == req_index | valid_31; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_558 = 8'h20 == req_index | valid_32; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_559 = 8'h21 == req_index | valid_33; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_560 = 8'h22 == req_index | valid_34; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_561 = 8'h23 == req_index | valid_35; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_562 = 8'h24 == req_index | valid_36; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_563 = 8'h25 == req_index | valid_37; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_564 = 8'h26 == req_index | valid_38; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_565 = 8'h27 == req_index | valid_39; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_566 = 8'h28 == req_index | valid_40; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_567 = 8'h29 == req_index | valid_41; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_568 = 8'h2a == req_index | valid_42; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_569 = 8'h2b == req_index | valid_43; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_570 = 8'h2c == req_index | valid_44; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_571 = 8'h2d == req_index | valid_45; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_572 = 8'h2e == req_index | valid_46; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_573 = 8'h2f == req_index | valid_47; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_574 = 8'h30 == req_index | valid_48; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_575 = 8'h31 == req_index | valid_49; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_576 = 8'h32 == req_index | valid_50; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_577 = 8'h33 == req_index | valid_51; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_578 = 8'h34 == req_index | valid_52; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_579 = 8'h35 == req_index | valid_53; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_580 = 8'h36 == req_index | valid_54; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_581 = 8'h37 == req_index | valid_55; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_582 = 8'h38 == req_index | valid_56; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_583 = 8'h39 == req_index | valid_57; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_584 = 8'h3a == req_index | valid_58; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_585 = 8'h3b == req_index | valid_59; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_586 = 8'h3c == req_index | valid_60; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_587 = 8'h3d == req_index | valid_61; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_588 = 8'h3e == req_index | valid_62; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_589 = 8'h3f == req_index | valid_63; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_590 = 8'h40 == req_index | valid_64; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_591 = 8'h41 == req_index | valid_65; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_592 = 8'h42 == req_index | valid_66; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_593 = 8'h43 == req_index | valid_67; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_594 = 8'h44 == req_index | valid_68; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_595 = 8'h45 == req_index | valid_69; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_596 = 8'h46 == req_index | valid_70; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_597 = 8'h47 == req_index | valid_71; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_598 = 8'h48 == req_index | valid_72; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_599 = 8'h49 == req_index | valid_73; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_600 = 8'h4a == req_index | valid_74; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_601 = 8'h4b == req_index | valid_75; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_602 = 8'h4c == req_index | valid_76; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_603 = 8'h4d == req_index | valid_77; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_604 = 8'h4e == req_index | valid_78; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_605 = 8'h4f == req_index | valid_79; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_606 = 8'h50 == req_index | valid_80; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_607 = 8'h51 == req_index | valid_81; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_608 = 8'h52 == req_index | valid_82; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_609 = 8'h53 == req_index | valid_83; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_610 = 8'h54 == req_index | valid_84; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_611 = 8'h55 == req_index | valid_85; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_612 = 8'h56 == req_index | valid_86; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_613 = 8'h57 == req_index | valid_87; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_614 = 8'h58 == req_index | valid_88; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_615 = 8'h59 == req_index | valid_89; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_616 = 8'h5a == req_index | valid_90; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_617 = 8'h5b == req_index | valid_91; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_618 = 8'h5c == req_index | valid_92; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_619 = 8'h5d == req_index | valid_93; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_620 = 8'h5e == req_index | valid_94; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_621 = 8'h5f == req_index | valid_95; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_622 = 8'h60 == req_index | valid_96; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_623 = 8'h61 == req_index | valid_97; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_624 = 8'h62 == req_index | valid_98; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_625 = 8'h63 == req_index | valid_99; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_626 = 8'h64 == req_index | valid_100; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_627 = 8'h65 == req_index | valid_101; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_628 = 8'h66 == req_index | valid_102; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_629 = 8'h67 == req_index | valid_103; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_630 = 8'h68 == req_index | valid_104; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_631 = 8'h69 == req_index | valid_105; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_632 = 8'h6a == req_index | valid_106; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_633 = 8'h6b == req_index | valid_107; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_634 = 8'h6c == req_index | valid_108; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_635 = 8'h6d == req_index | valid_109; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_636 = 8'h6e == req_index | valid_110; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_637 = 8'h6f == req_index | valid_111; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_638 = 8'h70 == req_index | valid_112; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_639 = 8'h71 == req_index | valid_113; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_640 = 8'h72 == req_index | valid_114; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_641 = 8'h73 == req_index | valid_115; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_642 = 8'h74 == req_index | valid_116; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_643 = 8'h75 == req_index | valid_117; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_644 = 8'h76 == req_index | valid_118; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_645 = 8'h77 == req_index | valid_119; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_646 = 8'h78 == req_index | valid_120; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_647 = 8'h79 == req_index | valid_121; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_648 = 8'h7a == req_index | valid_122; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_649 = 8'h7b == req_index | valid_123; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_650 = 8'h7c == req_index | valid_124; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_651 = 8'h7d == req_index | valid_125; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_652 = 8'h7e == req_index | valid_126; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_653 = 8'h7f == req_index | valid_127; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_654 = 8'h80 == req_index | valid_128; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_655 = 8'h81 == req_index | valid_129; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_656 = 8'h82 == req_index | valid_130; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_657 = 8'h83 == req_index | valid_131; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_658 = 8'h84 == req_index | valid_132; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_659 = 8'h85 == req_index | valid_133; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_660 = 8'h86 == req_index | valid_134; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_661 = 8'h87 == req_index | valid_135; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_662 = 8'h88 == req_index | valid_136; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_663 = 8'h89 == req_index | valid_137; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_664 = 8'h8a == req_index | valid_138; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_665 = 8'h8b == req_index | valid_139; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_666 = 8'h8c == req_index | valid_140; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_667 = 8'h8d == req_index | valid_141; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_668 = 8'h8e == req_index | valid_142; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_669 = 8'h8f == req_index | valid_143; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_670 = 8'h90 == req_index | valid_144; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_671 = 8'h91 == req_index | valid_145; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_672 = 8'h92 == req_index | valid_146; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_673 = 8'h93 == req_index | valid_147; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_674 = 8'h94 == req_index | valid_148; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_675 = 8'h95 == req_index | valid_149; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_676 = 8'h96 == req_index | valid_150; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_677 = 8'h97 == req_index | valid_151; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_678 = 8'h98 == req_index | valid_152; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_679 = 8'h99 == req_index | valid_153; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_680 = 8'h9a == req_index | valid_154; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_681 = 8'h9b == req_index | valid_155; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_682 = 8'h9c == req_index | valid_156; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_683 = 8'h9d == req_index | valid_157; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_684 = 8'h9e == req_index | valid_158; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_685 = 8'h9f == req_index | valid_159; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_686 = 8'ha0 == req_index | valid_160; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_687 = 8'ha1 == req_index | valid_161; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_688 = 8'ha2 == req_index | valid_162; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_689 = 8'ha3 == req_index | valid_163; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_690 = 8'ha4 == req_index | valid_164; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_691 = 8'ha5 == req_index | valid_165; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_692 = 8'ha6 == req_index | valid_166; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_693 = 8'ha7 == req_index | valid_167; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_694 = 8'ha8 == req_index | valid_168; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_695 = 8'ha9 == req_index | valid_169; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_696 = 8'haa == req_index | valid_170; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_697 = 8'hab == req_index | valid_171; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_698 = 8'hac == req_index | valid_172; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_699 = 8'had == req_index | valid_173; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_700 = 8'hae == req_index | valid_174; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_701 = 8'haf == req_index | valid_175; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_702 = 8'hb0 == req_index | valid_176; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_703 = 8'hb1 == req_index | valid_177; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_704 = 8'hb2 == req_index | valid_178; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_705 = 8'hb3 == req_index | valid_179; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_706 = 8'hb4 == req_index | valid_180; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_707 = 8'hb5 == req_index | valid_181; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_708 = 8'hb6 == req_index | valid_182; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_709 = 8'hb7 == req_index | valid_183; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_710 = 8'hb8 == req_index | valid_184; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_711 = 8'hb9 == req_index | valid_185; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_712 = 8'hba == req_index | valid_186; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_713 = 8'hbb == req_index | valid_187; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_714 = 8'hbc == req_index | valid_188; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_715 = 8'hbd == req_index | valid_189; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_716 = 8'hbe == req_index | valid_190; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_717 = 8'hbf == req_index | valid_191; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_718 = 8'hc0 == req_index | valid_192; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_719 = 8'hc1 == req_index | valid_193; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_720 = 8'hc2 == req_index | valid_194; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_721 = 8'hc3 == req_index | valid_195; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_722 = 8'hc4 == req_index | valid_196; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_723 = 8'hc5 == req_index | valid_197; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_724 = 8'hc6 == req_index | valid_198; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_725 = 8'hc7 == req_index | valid_199; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_726 = 8'hc8 == req_index | valid_200; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_727 = 8'hc9 == req_index | valid_201; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_728 = 8'hca == req_index | valid_202; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_729 = 8'hcb == req_index | valid_203; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_730 = 8'hcc == req_index | valid_204; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_731 = 8'hcd == req_index | valid_205; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_732 = 8'hce == req_index | valid_206; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_733 = 8'hcf == req_index | valid_207; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_734 = 8'hd0 == req_index | valid_208; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_735 = 8'hd1 == req_index | valid_209; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_736 = 8'hd2 == req_index | valid_210; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_737 = 8'hd3 == req_index | valid_211; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_738 = 8'hd4 == req_index | valid_212; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_739 = 8'hd5 == req_index | valid_213; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_740 = 8'hd6 == req_index | valid_214; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_741 = 8'hd7 == req_index | valid_215; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_742 = 8'hd8 == req_index | valid_216; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_743 = 8'hd9 == req_index | valid_217; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_744 = 8'hda == req_index | valid_218; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_745 = 8'hdb == req_index | valid_219; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_746 = 8'hdc == req_index | valid_220; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_747 = 8'hdd == req_index | valid_221; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_748 = 8'hde == req_index | valid_222; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_749 = 8'hdf == req_index | valid_223; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_750 = 8'he0 == req_index | valid_224; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_751 = 8'he1 == req_index | valid_225; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_752 = 8'he2 == req_index | valid_226; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_753 = 8'he3 == req_index | valid_227; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_754 = 8'he4 == req_index | valid_228; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_755 = 8'he5 == req_index | valid_229; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_756 = 8'he6 == req_index | valid_230; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_757 = 8'he7 == req_index | valid_231; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_758 = 8'he8 == req_index | valid_232; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_759 = 8'he9 == req_index | valid_233; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_760 = 8'hea == req_index | valid_234; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_761 = 8'heb == req_index | valid_235; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_762 = 8'hec == req_index | valid_236; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_763 = 8'hed == req_index | valid_237; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_764 = 8'hee == req_index | valid_238; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_765 = 8'hef == req_index | valid_239; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_766 = 8'hf0 == req_index | valid_240; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_767 = 8'hf1 == req_index | valid_241; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_768 = 8'hf2 == req_index | valid_242; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_769 = 8'hf3 == req_index | valid_243; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_770 = 8'hf4 == req_index | valid_244; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_771 = 8'hf5 == req_index | valid_245; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_772 = 8'hf6 == req_index | valid_246; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_773 = 8'hf7 == req_index | valid_247; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_774 = 8'hf8 == req_index | valid_248; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_775 = 8'hf9 == req_index | valid_249; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_776 = 8'hfa == req_index | valid_250; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_777 = 8'hfb == req_index | valid_251; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_778 = 8'hfc == req_index | valid_252; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_779 = 8'hfd == req_index | valid_253; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_780 = 8'hfe == req_index | valid_254; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire  _GEN_781 = 8'hff == req_index | valid_255; // @[Icache.scala 100:25 Icache.scala 100:25 Icache.scala 17:24]
  wire [19:0] _GEN_782 = 8'h0 == req_index ? req_tag : tag_0; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_783 = 8'h1 == req_index ? req_tag : tag_1; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_784 = 8'h2 == req_index ? req_tag : tag_2; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_785 = 8'h3 == req_index ? req_tag : tag_3; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_786 = 8'h4 == req_index ? req_tag : tag_4; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_787 = 8'h5 == req_index ? req_tag : tag_5; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_788 = 8'h6 == req_index ? req_tag : tag_6; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_789 = 8'h7 == req_index ? req_tag : tag_7; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_790 = 8'h8 == req_index ? req_tag : tag_8; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_791 = 8'h9 == req_index ? req_tag : tag_9; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_792 = 8'ha == req_index ? req_tag : tag_10; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_793 = 8'hb == req_index ? req_tag : tag_11; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_794 = 8'hc == req_index ? req_tag : tag_12; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_795 = 8'hd == req_index ? req_tag : tag_13; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_796 = 8'he == req_index ? req_tag : tag_14; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_797 = 8'hf == req_index ? req_tag : tag_15; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_798 = 8'h10 == req_index ? req_tag : tag_16; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_799 = 8'h11 == req_index ? req_tag : tag_17; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_800 = 8'h12 == req_index ? req_tag : tag_18; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_801 = 8'h13 == req_index ? req_tag : tag_19; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_802 = 8'h14 == req_index ? req_tag : tag_20; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_803 = 8'h15 == req_index ? req_tag : tag_21; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_804 = 8'h16 == req_index ? req_tag : tag_22; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_805 = 8'h17 == req_index ? req_tag : tag_23; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_806 = 8'h18 == req_index ? req_tag : tag_24; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_807 = 8'h19 == req_index ? req_tag : tag_25; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_808 = 8'h1a == req_index ? req_tag : tag_26; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_809 = 8'h1b == req_index ? req_tag : tag_27; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_810 = 8'h1c == req_index ? req_tag : tag_28; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_811 = 8'h1d == req_index ? req_tag : tag_29; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_812 = 8'h1e == req_index ? req_tag : tag_30; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_813 = 8'h1f == req_index ? req_tag : tag_31; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_814 = 8'h20 == req_index ? req_tag : tag_32; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_815 = 8'h21 == req_index ? req_tag : tag_33; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_816 = 8'h22 == req_index ? req_tag : tag_34; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_817 = 8'h23 == req_index ? req_tag : tag_35; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_818 = 8'h24 == req_index ? req_tag : tag_36; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_819 = 8'h25 == req_index ? req_tag : tag_37; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_820 = 8'h26 == req_index ? req_tag : tag_38; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_821 = 8'h27 == req_index ? req_tag : tag_39; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_822 = 8'h28 == req_index ? req_tag : tag_40; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_823 = 8'h29 == req_index ? req_tag : tag_41; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_824 = 8'h2a == req_index ? req_tag : tag_42; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_825 = 8'h2b == req_index ? req_tag : tag_43; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_826 = 8'h2c == req_index ? req_tag : tag_44; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_827 = 8'h2d == req_index ? req_tag : tag_45; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_828 = 8'h2e == req_index ? req_tag : tag_46; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_829 = 8'h2f == req_index ? req_tag : tag_47; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_830 = 8'h30 == req_index ? req_tag : tag_48; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_831 = 8'h31 == req_index ? req_tag : tag_49; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_832 = 8'h32 == req_index ? req_tag : tag_50; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_833 = 8'h33 == req_index ? req_tag : tag_51; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_834 = 8'h34 == req_index ? req_tag : tag_52; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_835 = 8'h35 == req_index ? req_tag : tag_53; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_836 = 8'h36 == req_index ? req_tag : tag_54; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_837 = 8'h37 == req_index ? req_tag : tag_55; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_838 = 8'h38 == req_index ? req_tag : tag_56; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_839 = 8'h39 == req_index ? req_tag : tag_57; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_840 = 8'h3a == req_index ? req_tag : tag_58; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_841 = 8'h3b == req_index ? req_tag : tag_59; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_842 = 8'h3c == req_index ? req_tag : tag_60; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_843 = 8'h3d == req_index ? req_tag : tag_61; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_844 = 8'h3e == req_index ? req_tag : tag_62; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_845 = 8'h3f == req_index ? req_tag : tag_63; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_846 = 8'h40 == req_index ? req_tag : tag_64; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_847 = 8'h41 == req_index ? req_tag : tag_65; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_848 = 8'h42 == req_index ? req_tag : tag_66; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_849 = 8'h43 == req_index ? req_tag : tag_67; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_850 = 8'h44 == req_index ? req_tag : tag_68; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_851 = 8'h45 == req_index ? req_tag : tag_69; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_852 = 8'h46 == req_index ? req_tag : tag_70; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_853 = 8'h47 == req_index ? req_tag : tag_71; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_854 = 8'h48 == req_index ? req_tag : tag_72; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_855 = 8'h49 == req_index ? req_tag : tag_73; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_856 = 8'h4a == req_index ? req_tag : tag_74; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_857 = 8'h4b == req_index ? req_tag : tag_75; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_858 = 8'h4c == req_index ? req_tag : tag_76; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_859 = 8'h4d == req_index ? req_tag : tag_77; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_860 = 8'h4e == req_index ? req_tag : tag_78; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_861 = 8'h4f == req_index ? req_tag : tag_79; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_862 = 8'h50 == req_index ? req_tag : tag_80; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_863 = 8'h51 == req_index ? req_tag : tag_81; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_864 = 8'h52 == req_index ? req_tag : tag_82; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_865 = 8'h53 == req_index ? req_tag : tag_83; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_866 = 8'h54 == req_index ? req_tag : tag_84; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_867 = 8'h55 == req_index ? req_tag : tag_85; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_868 = 8'h56 == req_index ? req_tag : tag_86; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_869 = 8'h57 == req_index ? req_tag : tag_87; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_870 = 8'h58 == req_index ? req_tag : tag_88; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_871 = 8'h59 == req_index ? req_tag : tag_89; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_872 = 8'h5a == req_index ? req_tag : tag_90; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_873 = 8'h5b == req_index ? req_tag : tag_91; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_874 = 8'h5c == req_index ? req_tag : tag_92; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_875 = 8'h5d == req_index ? req_tag : tag_93; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_876 = 8'h5e == req_index ? req_tag : tag_94; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_877 = 8'h5f == req_index ? req_tag : tag_95; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_878 = 8'h60 == req_index ? req_tag : tag_96; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_879 = 8'h61 == req_index ? req_tag : tag_97; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_880 = 8'h62 == req_index ? req_tag : tag_98; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_881 = 8'h63 == req_index ? req_tag : tag_99; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_882 = 8'h64 == req_index ? req_tag : tag_100; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_883 = 8'h65 == req_index ? req_tag : tag_101; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_884 = 8'h66 == req_index ? req_tag : tag_102; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_885 = 8'h67 == req_index ? req_tag : tag_103; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_886 = 8'h68 == req_index ? req_tag : tag_104; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_887 = 8'h69 == req_index ? req_tag : tag_105; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_888 = 8'h6a == req_index ? req_tag : tag_106; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_889 = 8'h6b == req_index ? req_tag : tag_107; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_890 = 8'h6c == req_index ? req_tag : tag_108; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_891 = 8'h6d == req_index ? req_tag : tag_109; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_892 = 8'h6e == req_index ? req_tag : tag_110; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_893 = 8'h6f == req_index ? req_tag : tag_111; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_894 = 8'h70 == req_index ? req_tag : tag_112; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_895 = 8'h71 == req_index ? req_tag : tag_113; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_896 = 8'h72 == req_index ? req_tag : tag_114; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_897 = 8'h73 == req_index ? req_tag : tag_115; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_898 = 8'h74 == req_index ? req_tag : tag_116; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_899 = 8'h75 == req_index ? req_tag : tag_117; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_900 = 8'h76 == req_index ? req_tag : tag_118; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_901 = 8'h77 == req_index ? req_tag : tag_119; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_902 = 8'h78 == req_index ? req_tag : tag_120; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_903 = 8'h79 == req_index ? req_tag : tag_121; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_904 = 8'h7a == req_index ? req_tag : tag_122; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_905 = 8'h7b == req_index ? req_tag : tag_123; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_906 = 8'h7c == req_index ? req_tag : tag_124; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_907 = 8'h7d == req_index ? req_tag : tag_125; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_908 = 8'h7e == req_index ? req_tag : tag_126; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_909 = 8'h7f == req_index ? req_tag : tag_127; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_910 = 8'h80 == req_index ? req_tag : tag_128; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_911 = 8'h81 == req_index ? req_tag : tag_129; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_912 = 8'h82 == req_index ? req_tag : tag_130; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_913 = 8'h83 == req_index ? req_tag : tag_131; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_914 = 8'h84 == req_index ? req_tag : tag_132; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_915 = 8'h85 == req_index ? req_tag : tag_133; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_916 = 8'h86 == req_index ? req_tag : tag_134; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_917 = 8'h87 == req_index ? req_tag : tag_135; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_918 = 8'h88 == req_index ? req_tag : tag_136; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_919 = 8'h89 == req_index ? req_tag : tag_137; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_920 = 8'h8a == req_index ? req_tag : tag_138; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_921 = 8'h8b == req_index ? req_tag : tag_139; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_922 = 8'h8c == req_index ? req_tag : tag_140; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_923 = 8'h8d == req_index ? req_tag : tag_141; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_924 = 8'h8e == req_index ? req_tag : tag_142; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_925 = 8'h8f == req_index ? req_tag : tag_143; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_926 = 8'h90 == req_index ? req_tag : tag_144; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_927 = 8'h91 == req_index ? req_tag : tag_145; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_928 = 8'h92 == req_index ? req_tag : tag_146; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_929 = 8'h93 == req_index ? req_tag : tag_147; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_930 = 8'h94 == req_index ? req_tag : tag_148; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_931 = 8'h95 == req_index ? req_tag : tag_149; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_932 = 8'h96 == req_index ? req_tag : tag_150; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_933 = 8'h97 == req_index ? req_tag : tag_151; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_934 = 8'h98 == req_index ? req_tag : tag_152; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_935 = 8'h99 == req_index ? req_tag : tag_153; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_936 = 8'h9a == req_index ? req_tag : tag_154; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_937 = 8'h9b == req_index ? req_tag : tag_155; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_938 = 8'h9c == req_index ? req_tag : tag_156; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_939 = 8'h9d == req_index ? req_tag : tag_157; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_940 = 8'h9e == req_index ? req_tag : tag_158; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_941 = 8'h9f == req_index ? req_tag : tag_159; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_942 = 8'ha0 == req_index ? req_tag : tag_160; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_943 = 8'ha1 == req_index ? req_tag : tag_161; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_944 = 8'ha2 == req_index ? req_tag : tag_162; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_945 = 8'ha3 == req_index ? req_tag : tag_163; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_946 = 8'ha4 == req_index ? req_tag : tag_164; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_947 = 8'ha5 == req_index ? req_tag : tag_165; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_948 = 8'ha6 == req_index ? req_tag : tag_166; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_949 = 8'ha7 == req_index ? req_tag : tag_167; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_950 = 8'ha8 == req_index ? req_tag : tag_168; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_951 = 8'ha9 == req_index ? req_tag : tag_169; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_952 = 8'haa == req_index ? req_tag : tag_170; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_953 = 8'hab == req_index ? req_tag : tag_171; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_954 = 8'hac == req_index ? req_tag : tag_172; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_955 = 8'had == req_index ? req_tag : tag_173; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_956 = 8'hae == req_index ? req_tag : tag_174; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_957 = 8'haf == req_index ? req_tag : tag_175; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_958 = 8'hb0 == req_index ? req_tag : tag_176; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_959 = 8'hb1 == req_index ? req_tag : tag_177; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_960 = 8'hb2 == req_index ? req_tag : tag_178; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_961 = 8'hb3 == req_index ? req_tag : tag_179; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_962 = 8'hb4 == req_index ? req_tag : tag_180; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_963 = 8'hb5 == req_index ? req_tag : tag_181; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_964 = 8'hb6 == req_index ? req_tag : tag_182; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_965 = 8'hb7 == req_index ? req_tag : tag_183; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_966 = 8'hb8 == req_index ? req_tag : tag_184; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_967 = 8'hb9 == req_index ? req_tag : tag_185; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_968 = 8'hba == req_index ? req_tag : tag_186; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_969 = 8'hbb == req_index ? req_tag : tag_187; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_970 = 8'hbc == req_index ? req_tag : tag_188; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_971 = 8'hbd == req_index ? req_tag : tag_189; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_972 = 8'hbe == req_index ? req_tag : tag_190; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_973 = 8'hbf == req_index ? req_tag : tag_191; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_974 = 8'hc0 == req_index ? req_tag : tag_192; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_975 = 8'hc1 == req_index ? req_tag : tag_193; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_976 = 8'hc2 == req_index ? req_tag : tag_194; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_977 = 8'hc3 == req_index ? req_tag : tag_195; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_978 = 8'hc4 == req_index ? req_tag : tag_196; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_979 = 8'hc5 == req_index ? req_tag : tag_197; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_980 = 8'hc6 == req_index ? req_tag : tag_198; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_981 = 8'hc7 == req_index ? req_tag : tag_199; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_982 = 8'hc8 == req_index ? req_tag : tag_200; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_983 = 8'hc9 == req_index ? req_tag : tag_201; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_984 = 8'hca == req_index ? req_tag : tag_202; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_985 = 8'hcb == req_index ? req_tag : tag_203; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_986 = 8'hcc == req_index ? req_tag : tag_204; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_987 = 8'hcd == req_index ? req_tag : tag_205; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_988 = 8'hce == req_index ? req_tag : tag_206; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_989 = 8'hcf == req_index ? req_tag : tag_207; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_990 = 8'hd0 == req_index ? req_tag : tag_208; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_991 = 8'hd1 == req_index ? req_tag : tag_209; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_992 = 8'hd2 == req_index ? req_tag : tag_210; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_993 = 8'hd3 == req_index ? req_tag : tag_211; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_994 = 8'hd4 == req_index ? req_tag : tag_212; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_995 = 8'hd5 == req_index ? req_tag : tag_213; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_996 = 8'hd6 == req_index ? req_tag : tag_214; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_997 = 8'hd7 == req_index ? req_tag : tag_215; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_998 = 8'hd8 == req_index ? req_tag : tag_216; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_999 = 8'hd9 == req_index ? req_tag : tag_217; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1000 = 8'hda == req_index ? req_tag : tag_218; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1001 = 8'hdb == req_index ? req_tag : tag_219; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1002 = 8'hdc == req_index ? req_tag : tag_220; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1003 = 8'hdd == req_index ? req_tag : tag_221; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1004 = 8'hde == req_index ? req_tag : tag_222; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1005 = 8'hdf == req_index ? req_tag : tag_223; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1006 = 8'he0 == req_index ? req_tag : tag_224; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1007 = 8'he1 == req_index ? req_tag : tag_225; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1008 = 8'he2 == req_index ? req_tag : tag_226; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1009 = 8'he3 == req_index ? req_tag : tag_227; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1010 = 8'he4 == req_index ? req_tag : tag_228; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1011 = 8'he5 == req_index ? req_tag : tag_229; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1012 = 8'he6 == req_index ? req_tag : tag_230; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1013 = 8'he7 == req_index ? req_tag : tag_231; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1014 = 8'he8 == req_index ? req_tag : tag_232; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1015 = 8'he9 == req_index ? req_tag : tag_233; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1016 = 8'hea == req_index ? req_tag : tag_234; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1017 = 8'heb == req_index ? req_tag : tag_235; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1018 = 8'hec == req_index ? req_tag : tag_236; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1019 = 8'hed == req_index ? req_tag : tag_237; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1020 = 8'hee == req_index ? req_tag : tag_238; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1021 = 8'hef == req_index ? req_tag : tag_239; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1022 = 8'hf0 == req_index ? req_tag : tag_240; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1023 = 8'hf1 == req_index ? req_tag : tag_241; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1024 = 8'hf2 == req_index ? req_tag : tag_242; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1025 = 8'hf3 == req_index ? req_tag : tag_243; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1026 = 8'hf4 == req_index ? req_tag : tag_244; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1027 = 8'hf5 == req_index ? req_tag : tag_245; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1028 = 8'hf6 == req_index ? req_tag : tag_246; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1029 = 8'hf7 == req_index ? req_tag : tag_247; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1030 = 8'hf8 == req_index ? req_tag : tag_248; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1031 = 8'hf9 == req_index ? req_tag : tag_249; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1032 = 8'hfa == req_index ? req_tag : tag_250; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1033 = 8'hfb == req_index ? req_tag : tag_251; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1034 = 8'hfc == req_index ? req_tag : tag_252; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1035 = 8'hfd == req_index ? req_tag : tag_253; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1036 = 8'hfe == req_index ? req_tag : tag_254; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire [19:0] _GEN_1037 = 8'hff == req_index ? req_tag : tag_255; // @[Icache.scala 101:25 Icache.scala 101:25 Icache.scala 16:24]
  wire  _GEN_1294 = _T_4 ? 1'h0 : cache_fill; // @[Conditional.scala 39:67 Icache.scala 98:25 Icache.scala 51:28]
  wire  _GEN_1295 = _T_4 ? 1'h0 : cache_wen; // @[Conditional.scala 39:67 Icache.scala 99:25 Icache.scala 52:28]
  wire  _GEN_1296 = _T_4 ? _GEN_526 : valid_0; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1297 = _T_4 ? _GEN_527 : valid_1; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1298 = _T_4 ? _GEN_528 : valid_2; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1299 = _T_4 ? _GEN_529 : valid_3; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1300 = _T_4 ? _GEN_530 : valid_4; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1301 = _T_4 ? _GEN_531 : valid_5; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1302 = _T_4 ? _GEN_532 : valid_6; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1303 = _T_4 ? _GEN_533 : valid_7; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1304 = _T_4 ? _GEN_534 : valid_8; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1305 = _T_4 ? _GEN_535 : valid_9; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1306 = _T_4 ? _GEN_536 : valid_10; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1307 = _T_4 ? _GEN_537 : valid_11; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1308 = _T_4 ? _GEN_538 : valid_12; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1309 = _T_4 ? _GEN_539 : valid_13; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1310 = _T_4 ? _GEN_540 : valid_14; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1311 = _T_4 ? _GEN_541 : valid_15; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1312 = _T_4 ? _GEN_542 : valid_16; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1313 = _T_4 ? _GEN_543 : valid_17; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1314 = _T_4 ? _GEN_544 : valid_18; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1315 = _T_4 ? _GEN_545 : valid_19; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1316 = _T_4 ? _GEN_546 : valid_20; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1317 = _T_4 ? _GEN_547 : valid_21; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1318 = _T_4 ? _GEN_548 : valid_22; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1319 = _T_4 ? _GEN_549 : valid_23; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1320 = _T_4 ? _GEN_550 : valid_24; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1321 = _T_4 ? _GEN_551 : valid_25; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1322 = _T_4 ? _GEN_552 : valid_26; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1323 = _T_4 ? _GEN_553 : valid_27; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1324 = _T_4 ? _GEN_554 : valid_28; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1325 = _T_4 ? _GEN_555 : valid_29; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1326 = _T_4 ? _GEN_556 : valid_30; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1327 = _T_4 ? _GEN_557 : valid_31; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1328 = _T_4 ? _GEN_558 : valid_32; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1329 = _T_4 ? _GEN_559 : valid_33; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1330 = _T_4 ? _GEN_560 : valid_34; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1331 = _T_4 ? _GEN_561 : valid_35; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1332 = _T_4 ? _GEN_562 : valid_36; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1333 = _T_4 ? _GEN_563 : valid_37; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1334 = _T_4 ? _GEN_564 : valid_38; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1335 = _T_4 ? _GEN_565 : valid_39; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1336 = _T_4 ? _GEN_566 : valid_40; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1337 = _T_4 ? _GEN_567 : valid_41; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1338 = _T_4 ? _GEN_568 : valid_42; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1339 = _T_4 ? _GEN_569 : valid_43; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1340 = _T_4 ? _GEN_570 : valid_44; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1341 = _T_4 ? _GEN_571 : valid_45; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1342 = _T_4 ? _GEN_572 : valid_46; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1343 = _T_4 ? _GEN_573 : valid_47; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1344 = _T_4 ? _GEN_574 : valid_48; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1345 = _T_4 ? _GEN_575 : valid_49; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1346 = _T_4 ? _GEN_576 : valid_50; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1347 = _T_4 ? _GEN_577 : valid_51; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1348 = _T_4 ? _GEN_578 : valid_52; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1349 = _T_4 ? _GEN_579 : valid_53; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1350 = _T_4 ? _GEN_580 : valid_54; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1351 = _T_4 ? _GEN_581 : valid_55; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1352 = _T_4 ? _GEN_582 : valid_56; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1353 = _T_4 ? _GEN_583 : valid_57; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1354 = _T_4 ? _GEN_584 : valid_58; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1355 = _T_4 ? _GEN_585 : valid_59; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1356 = _T_4 ? _GEN_586 : valid_60; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1357 = _T_4 ? _GEN_587 : valid_61; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1358 = _T_4 ? _GEN_588 : valid_62; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1359 = _T_4 ? _GEN_589 : valid_63; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1360 = _T_4 ? _GEN_590 : valid_64; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1361 = _T_4 ? _GEN_591 : valid_65; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1362 = _T_4 ? _GEN_592 : valid_66; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1363 = _T_4 ? _GEN_593 : valid_67; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1364 = _T_4 ? _GEN_594 : valid_68; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1365 = _T_4 ? _GEN_595 : valid_69; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1366 = _T_4 ? _GEN_596 : valid_70; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1367 = _T_4 ? _GEN_597 : valid_71; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1368 = _T_4 ? _GEN_598 : valid_72; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1369 = _T_4 ? _GEN_599 : valid_73; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1370 = _T_4 ? _GEN_600 : valid_74; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1371 = _T_4 ? _GEN_601 : valid_75; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1372 = _T_4 ? _GEN_602 : valid_76; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1373 = _T_4 ? _GEN_603 : valid_77; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1374 = _T_4 ? _GEN_604 : valid_78; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1375 = _T_4 ? _GEN_605 : valid_79; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1376 = _T_4 ? _GEN_606 : valid_80; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1377 = _T_4 ? _GEN_607 : valid_81; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1378 = _T_4 ? _GEN_608 : valid_82; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1379 = _T_4 ? _GEN_609 : valid_83; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1380 = _T_4 ? _GEN_610 : valid_84; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1381 = _T_4 ? _GEN_611 : valid_85; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1382 = _T_4 ? _GEN_612 : valid_86; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1383 = _T_4 ? _GEN_613 : valid_87; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1384 = _T_4 ? _GEN_614 : valid_88; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1385 = _T_4 ? _GEN_615 : valid_89; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1386 = _T_4 ? _GEN_616 : valid_90; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1387 = _T_4 ? _GEN_617 : valid_91; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1388 = _T_4 ? _GEN_618 : valid_92; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1389 = _T_4 ? _GEN_619 : valid_93; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1390 = _T_4 ? _GEN_620 : valid_94; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1391 = _T_4 ? _GEN_621 : valid_95; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1392 = _T_4 ? _GEN_622 : valid_96; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1393 = _T_4 ? _GEN_623 : valid_97; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1394 = _T_4 ? _GEN_624 : valid_98; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1395 = _T_4 ? _GEN_625 : valid_99; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1396 = _T_4 ? _GEN_626 : valid_100; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1397 = _T_4 ? _GEN_627 : valid_101; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1398 = _T_4 ? _GEN_628 : valid_102; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1399 = _T_4 ? _GEN_629 : valid_103; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1400 = _T_4 ? _GEN_630 : valid_104; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1401 = _T_4 ? _GEN_631 : valid_105; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1402 = _T_4 ? _GEN_632 : valid_106; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1403 = _T_4 ? _GEN_633 : valid_107; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1404 = _T_4 ? _GEN_634 : valid_108; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1405 = _T_4 ? _GEN_635 : valid_109; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1406 = _T_4 ? _GEN_636 : valid_110; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1407 = _T_4 ? _GEN_637 : valid_111; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1408 = _T_4 ? _GEN_638 : valid_112; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1409 = _T_4 ? _GEN_639 : valid_113; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1410 = _T_4 ? _GEN_640 : valid_114; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1411 = _T_4 ? _GEN_641 : valid_115; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1412 = _T_4 ? _GEN_642 : valid_116; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1413 = _T_4 ? _GEN_643 : valid_117; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1414 = _T_4 ? _GEN_644 : valid_118; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1415 = _T_4 ? _GEN_645 : valid_119; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1416 = _T_4 ? _GEN_646 : valid_120; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1417 = _T_4 ? _GEN_647 : valid_121; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1418 = _T_4 ? _GEN_648 : valid_122; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1419 = _T_4 ? _GEN_649 : valid_123; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1420 = _T_4 ? _GEN_650 : valid_124; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1421 = _T_4 ? _GEN_651 : valid_125; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1422 = _T_4 ? _GEN_652 : valid_126; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1423 = _T_4 ? _GEN_653 : valid_127; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1424 = _T_4 ? _GEN_654 : valid_128; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1425 = _T_4 ? _GEN_655 : valid_129; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1426 = _T_4 ? _GEN_656 : valid_130; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1427 = _T_4 ? _GEN_657 : valid_131; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1428 = _T_4 ? _GEN_658 : valid_132; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1429 = _T_4 ? _GEN_659 : valid_133; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1430 = _T_4 ? _GEN_660 : valid_134; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1431 = _T_4 ? _GEN_661 : valid_135; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1432 = _T_4 ? _GEN_662 : valid_136; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1433 = _T_4 ? _GEN_663 : valid_137; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1434 = _T_4 ? _GEN_664 : valid_138; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1435 = _T_4 ? _GEN_665 : valid_139; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1436 = _T_4 ? _GEN_666 : valid_140; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1437 = _T_4 ? _GEN_667 : valid_141; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1438 = _T_4 ? _GEN_668 : valid_142; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1439 = _T_4 ? _GEN_669 : valid_143; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1440 = _T_4 ? _GEN_670 : valid_144; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1441 = _T_4 ? _GEN_671 : valid_145; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1442 = _T_4 ? _GEN_672 : valid_146; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1443 = _T_4 ? _GEN_673 : valid_147; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1444 = _T_4 ? _GEN_674 : valid_148; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1445 = _T_4 ? _GEN_675 : valid_149; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1446 = _T_4 ? _GEN_676 : valid_150; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1447 = _T_4 ? _GEN_677 : valid_151; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1448 = _T_4 ? _GEN_678 : valid_152; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1449 = _T_4 ? _GEN_679 : valid_153; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1450 = _T_4 ? _GEN_680 : valid_154; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1451 = _T_4 ? _GEN_681 : valid_155; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1452 = _T_4 ? _GEN_682 : valid_156; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1453 = _T_4 ? _GEN_683 : valid_157; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1454 = _T_4 ? _GEN_684 : valid_158; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1455 = _T_4 ? _GEN_685 : valid_159; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1456 = _T_4 ? _GEN_686 : valid_160; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1457 = _T_4 ? _GEN_687 : valid_161; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1458 = _T_4 ? _GEN_688 : valid_162; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1459 = _T_4 ? _GEN_689 : valid_163; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1460 = _T_4 ? _GEN_690 : valid_164; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1461 = _T_4 ? _GEN_691 : valid_165; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1462 = _T_4 ? _GEN_692 : valid_166; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1463 = _T_4 ? _GEN_693 : valid_167; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1464 = _T_4 ? _GEN_694 : valid_168; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1465 = _T_4 ? _GEN_695 : valid_169; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1466 = _T_4 ? _GEN_696 : valid_170; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1467 = _T_4 ? _GEN_697 : valid_171; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1468 = _T_4 ? _GEN_698 : valid_172; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1469 = _T_4 ? _GEN_699 : valid_173; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1470 = _T_4 ? _GEN_700 : valid_174; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1471 = _T_4 ? _GEN_701 : valid_175; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1472 = _T_4 ? _GEN_702 : valid_176; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1473 = _T_4 ? _GEN_703 : valid_177; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1474 = _T_4 ? _GEN_704 : valid_178; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1475 = _T_4 ? _GEN_705 : valid_179; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1476 = _T_4 ? _GEN_706 : valid_180; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1477 = _T_4 ? _GEN_707 : valid_181; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1478 = _T_4 ? _GEN_708 : valid_182; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1479 = _T_4 ? _GEN_709 : valid_183; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1480 = _T_4 ? _GEN_710 : valid_184; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1481 = _T_4 ? _GEN_711 : valid_185; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1482 = _T_4 ? _GEN_712 : valid_186; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1483 = _T_4 ? _GEN_713 : valid_187; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1484 = _T_4 ? _GEN_714 : valid_188; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1485 = _T_4 ? _GEN_715 : valid_189; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1486 = _T_4 ? _GEN_716 : valid_190; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1487 = _T_4 ? _GEN_717 : valid_191; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1488 = _T_4 ? _GEN_718 : valid_192; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1489 = _T_4 ? _GEN_719 : valid_193; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1490 = _T_4 ? _GEN_720 : valid_194; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1491 = _T_4 ? _GEN_721 : valid_195; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1492 = _T_4 ? _GEN_722 : valid_196; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1493 = _T_4 ? _GEN_723 : valid_197; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1494 = _T_4 ? _GEN_724 : valid_198; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1495 = _T_4 ? _GEN_725 : valid_199; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1496 = _T_4 ? _GEN_726 : valid_200; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1497 = _T_4 ? _GEN_727 : valid_201; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1498 = _T_4 ? _GEN_728 : valid_202; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1499 = _T_4 ? _GEN_729 : valid_203; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1500 = _T_4 ? _GEN_730 : valid_204; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1501 = _T_4 ? _GEN_731 : valid_205; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1502 = _T_4 ? _GEN_732 : valid_206; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1503 = _T_4 ? _GEN_733 : valid_207; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1504 = _T_4 ? _GEN_734 : valid_208; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1505 = _T_4 ? _GEN_735 : valid_209; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1506 = _T_4 ? _GEN_736 : valid_210; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1507 = _T_4 ? _GEN_737 : valid_211; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1508 = _T_4 ? _GEN_738 : valid_212; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1509 = _T_4 ? _GEN_739 : valid_213; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1510 = _T_4 ? _GEN_740 : valid_214; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1511 = _T_4 ? _GEN_741 : valid_215; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1512 = _T_4 ? _GEN_742 : valid_216; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1513 = _T_4 ? _GEN_743 : valid_217; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1514 = _T_4 ? _GEN_744 : valid_218; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1515 = _T_4 ? _GEN_745 : valid_219; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1516 = _T_4 ? _GEN_746 : valid_220; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1517 = _T_4 ? _GEN_747 : valid_221; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1518 = _T_4 ? _GEN_748 : valid_222; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1519 = _T_4 ? _GEN_749 : valid_223; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1520 = _T_4 ? _GEN_750 : valid_224; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1521 = _T_4 ? _GEN_751 : valid_225; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1522 = _T_4 ? _GEN_752 : valid_226; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1523 = _T_4 ? _GEN_753 : valid_227; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1524 = _T_4 ? _GEN_754 : valid_228; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1525 = _T_4 ? _GEN_755 : valid_229; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1526 = _T_4 ? _GEN_756 : valid_230; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1527 = _T_4 ? _GEN_757 : valid_231; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1528 = _T_4 ? _GEN_758 : valid_232; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1529 = _T_4 ? _GEN_759 : valid_233; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1530 = _T_4 ? _GEN_760 : valid_234; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1531 = _T_4 ? _GEN_761 : valid_235; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1532 = _T_4 ? _GEN_762 : valid_236; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1533 = _T_4 ? _GEN_763 : valid_237; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1534 = _T_4 ? _GEN_764 : valid_238; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1535 = _T_4 ? _GEN_765 : valid_239; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1536 = _T_4 ? _GEN_766 : valid_240; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1537 = _T_4 ? _GEN_767 : valid_241; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1538 = _T_4 ? _GEN_768 : valid_242; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1539 = _T_4 ? _GEN_769 : valid_243; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1540 = _T_4 ? _GEN_770 : valid_244; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1541 = _T_4 ? _GEN_771 : valid_245; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1542 = _T_4 ? _GEN_772 : valid_246; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1543 = _T_4 ? _GEN_773 : valid_247; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1544 = _T_4 ? _GEN_774 : valid_248; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1545 = _T_4 ? _GEN_775 : valid_249; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1546 = _T_4 ? _GEN_776 : valid_250; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1547 = _T_4 ? _GEN_777 : valid_251; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1548 = _T_4 ? _GEN_778 : valid_252; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1549 = _T_4 ? _GEN_779 : valid_253; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1550 = _T_4 ? _GEN_780 : valid_254; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire  _GEN_1551 = _T_4 ? _GEN_781 : valid_255; // @[Conditional.scala 39:67 Icache.scala 17:24]
  wire [19:0] _GEN_1552 = _T_4 ? _GEN_782 : tag_0; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1553 = _T_4 ? _GEN_783 : tag_1; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1554 = _T_4 ? _GEN_784 : tag_2; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1555 = _T_4 ? _GEN_785 : tag_3; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1556 = _T_4 ? _GEN_786 : tag_4; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1557 = _T_4 ? _GEN_787 : tag_5; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1558 = _T_4 ? _GEN_788 : tag_6; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1559 = _T_4 ? _GEN_789 : tag_7; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1560 = _T_4 ? _GEN_790 : tag_8; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1561 = _T_4 ? _GEN_791 : tag_9; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1562 = _T_4 ? _GEN_792 : tag_10; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1563 = _T_4 ? _GEN_793 : tag_11; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1564 = _T_4 ? _GEN_794 : tag_12; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1565 = _T_4 ? _GEN_795 : tag_13; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1566 = _T_4 ? _GEN_796 : tag_14; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1567 = _T_4 ? _GEN_797 : tag_15; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1568 = _T_4 ? _GEN_798 : tag_16; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1569 = _T_4 ? _GEN_799 : tag_17; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1570 = _T_4 ? _GEN_800 : tag_18; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1571 = _T_4 ? _GEN_801 : tag_19; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1572 = _T_4 ? _GEN_802 : tag_20; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1573 = _T_4 ? _GEN_803 : tag_21; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1574 = _T_4 ? _GEN_804 : tag_22; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1575 = _T_4 ? _GEN_805 : tag_23; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1576 = _T_4 ? _GEN_806 : tag_24; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1577 = _T_4 ? _GEN_807 : tag_25; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1578 = _T_4 ? _GEN_808 : tag_26; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1579 = _T_4 ? _GEN_809 : tag_27; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1580 = _T_4 ? _GEN_810 : tag_28; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1581 = _T_4 ? _GEN_811 : tag_29; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1582 = _T_4 ? _GEN_812 : tag_30; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1583 = _T_4 ? _GEN_813 : tag_31; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1584 = _T_4 ? _GEN_814 : tag_32; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1585 = _T_4 ? _GEN_815 : tag_33; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1586 = _T_4 ? _GEN_816 : tag_34; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1587 = _T_4 ? _GEN_817 : tag_35; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1588 = _T_4 ? _GEN_818 : tag_36; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1589 = _T_4 ? _GEN_819 : tag_37; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1590 = _T_4 ? _GEN_820 : tag_38; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1591 = _T_4 ? _GEN_821 : tag_39; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1592 = _T_4 ? _GEN_822 : tag_40; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1593 = _T_4 ? _GEN_823 : tag_41; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1594 = _T_4 ? _GEN_824 : tag_42; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1595 = _T_4 ? _GEN_825 : tag_43; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1596 = _T_4 ? _GEN_826 : tag_44; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1597 = _T_4 ? _GEN_827 : tag_45; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1598 = _T_4 ? _GEN_828 : tag_46; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1599 = _T_4 ? _GEN_829 : tag_47; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1600 = _T_4 ? _GEN_830 : tag_48; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1601 = _T_4 ? _GEN_831 : tag_49; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1602 = _T_4 ? _GEN_832 : tag_50; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1603 = _T_4 ? _GEN_833 : tag_51; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1604 = _T_4 ? _GEN_834 : tag_52; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1605 = _T_4 ? _GEN_835 : tag_53; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1606 = _T_4 ? _GEN_836 : tag_54; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1607 = _T_4 ? _GEN_837 : tag_55; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1608 = _T_4 ? _GEN_838 : tag_56; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1609 = _T_4 ? _GEN_839 : tag_57; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1610 = _T_4 ? _GEN_840 : tag_58; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1611 = _T_4 ? _GEN_841 : tag_59; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1612 = _T_4 ? _GEN_842 : tag_60; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1613 = _T_4 ? _GEN_843 : tag_61; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1614 = _T_4 ? _GEN_844 : tag_62; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1615 = _T_4 ? _GEN_845 : tag_63; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1616 = _T_4 ? _GEN_846 : tag_64; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1617 = _T_4 ? _GEN_847 : tag_65; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1618 = _T_4 ? _GEN_848 : tag_66; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1619 = _T_4 ? _GEN_849 : tag_67; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1620 = _T_4 ? _GEN_850 : tag_68; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1621 = _T_4 ? _GEN_851 : tag_69; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1622 = _T_4 ? _GEN_852 : tag_70; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1623 = _T_4 ? _GEN_853 : tag_71; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1624 = _T_4 ? _GEN_854 : tag_72; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1625 = _T_4 ? _GEN_855 : tag_73; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1626 = _T_4 ? _GEN_856 : tag_74; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1627 = _T_4 ? _GEN_857 : tag_75; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1628 = _T_4 ? _GEN_858 : tag_76; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1629 = _T_4 ? _GEN_859 : tag_77; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1630 = _T_4 ? _GEN_860 : tag_78; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1631 = _T_4 ? _GEN_861 : tag_79; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1632 = _T_4 ? _GEN_862 : tag_80; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1633 = _T_4 ? _GEN_863 : tag_81; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1634 = _T_4 ? _GEN_864 : tag_82; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1635 = _T_4 ? _GEN_865 : tag_83; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1636 = _T_4 ? _GEN_866 : tag_84; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1637 = _T_4 ? _GEN_867 : tag_85; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1638 = _T_4 ? _GEN_868 : tag_86; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1639 = _T_4 ? _GEN_869 : tag_87; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1640 = _T_4 ? _GEN_870 : tag_88; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1641 = _T_4 ? _GEN_871 : tag_89; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1642 = _T_4 ? _GEN_872 : tag_90; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1643 = _T_4 ? _GEN_873 : tag_91; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1644 = _T_4 ? _GEN_874 : tag_92; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1645 = _T_4 ? _GEN_875 : tag_93; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1646 = _T_4 ? _GEN_876 : tag_94; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1647 = _T_4 ? _GEN_877 : tag_95; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1648 = _T_4 ? _GEN_878 : tag_96; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1649 = _T_4 ? _GEN_879 : tag_97; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1650 = _T_4 ? _GEN_880 : tag_98; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1651 = _T_4 ? _GEN_881 : tag_99; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1652 = _T_4 ? _GEN_882 : tag_100; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1653 = _T_4 ? _GEN_883 : tag_101; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1654 = _T_4 ? _GEN_884 : tag_102; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1655 = _T_4 ? _GEN_885 : tag_103; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1656 = _T_4 ? _GEN_886 : tag_104; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1657 = _T_4 ? _GEN_887 : tag_105; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1658 = _T_4 ? _GEN_888 : tag_106; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1659 = _T_4 ? _GEN_889 : tag_107; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1660 = _T_4 ? _GEN_890 : tag_108; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1661 = _T_4 ? _GEN_891 : tag_109; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1662 = _T_4 ? _GEN_892 : tag_110; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1663 = _T_4 ? _GEN_893 : tag_111; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1664 = _T_4 ? _GEN_894 : tag_112; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1665 = _T_4 ? _GEN_895 : tag_113; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1666 = _T_4 ? _GEN_896 : tag_114; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1667 = _T_4 ? _GEN_897 : tag_115; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1668 = _T_4 ? _GEN_898 : tag_116; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1669 = _T_4 ? _GEN_899 : tag_117; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1670 = _T_4 ? _GEN_900 : tag_118; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1671 = _T_4 ? _GEN_901 : tag_119; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1672 = _T_4 ? _GEN_902 : tag_120; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1673 = _T_4 ? _GEN_903 : tag_121; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1674 = _T_4 ? _GEN_904 : tag_122; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1675 = _T_4 ? _GEN_905 : tag_123; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1676 = _T_4 ? _GEN_906 : tag_124; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1677 = _T_4 ? _GEN_907 : tag_125; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1678 = _T_4 ? _GEN_908 : tag_126; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1679 = _T_4 ? _GEN_909 : tag_127; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1680 = _T_4 ? _GEN_910 : tag_128; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1681 = _T_4 ? _GEN_911 : tag_129; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1682 = _T_4 ? _GEN_912 : tag_130; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1683 = _T_4 ? _GEN_913 : tag_131; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1684 = _T_4 ? _GEN_914 : tag_132; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1685 = _T_4 ? _GEN_915 : tag_133; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1686 = _T_4 ? _GEN_916 : tag_134; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1687 = _T_4 ? _GEN_917 : tag_135; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1688 = _T_4 ? _GEN_918 : tag_136; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1689 = _T_4 ? _GEN_919 : tag_137; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1690 = _T_4 ? _GEN_920 : tag_138; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1691 = _T_4 ? _GEN_921 : tag_139; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1692 = _T_4 ? _GEN_922 : tag_140; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1693 = _T_4 ? _GEN_923 : tag_141; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1694 = _T_4 ? _GEN_924 : tag_142; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1695 = _T_4 ? _GEN_925 : tag_143; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1696 = _T_4 ? _GEN_926 : tag_144; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1697 = _T_4 ? _GEN_927 : tag_145; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1698 = _T_4 ? _GEN_928 : tag_146; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1699 = _T_4 ? _GEN_929 : tag_147; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1700 = _T_4 ? _GEN_930 : tag_148; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1701 = _T_4 ? _GEN_931 : tag_149; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1702 = _T_4 ? _GEN_932 : tag_150; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1703 = _T_4 ? _GEN_933 : tag_151; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1704 = _T_4 ? _GEN_934 : tag_152; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1705 = _T_4 ? _GEN_935 : tag_153; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1706 = _T_4 ? _GEN_936 : tag_154; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1707 = _T_4 ? _GEN_937 : tag_155; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1708 = _T_4 ? _GEN_938 : tag_156; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1709 = _T_4 ? _GEN_939 : tag_157; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1710 = _T_4 ? _GEN_940 : tag_158; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1711 = _T_4 ? _GEN_941 : tag_159; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1712 = _T_4 ? _GEN_942 : tag_160; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1713 = _T_4 ? _GEN_943 : tag_161; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1714 = _T_4 ? _GEN_944 : tag_162; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1715 = _T_4 ? _GEN_945 : tag_163; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1716 = _T_4 ? _GEN_946 : tag_164; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1717 = _T_4 ? _GEN_947 : tag_165; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1718 = _T_4 ? _GEN_948 : tag_166; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1719 = _T_4 ? _GEN_949 : tag_167; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1720 = _T_4 ? _GEN_950 : tag_168; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1721 = _T_4 ? _GEN_951 : tag_169; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1722 = _T_4 ? _GEN_952 : tag_170; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1723 = _T_4 ? _GEN_953 : tag_171; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1724 = _T_4 ? _GEN_954 : tag_172; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1725 = _T_4 ? _GEN_955 : tag_173; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1726 = _T_4 ? _GEN_956 : tag_174; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1727 = _T_4 ? _GEN_957 : tag_175; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1728 = _T_4 ? _GEN_958 : tag_176; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1729 = _T_4 ? _GEN_959 : tag_177; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1730 = _T_4 ? _GEN_960 : tag_178; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1731 = _T_4 ? _GEN_961 : tag_179; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1732 = _T_4 ? _GEN_962 : tag_180; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1733 = _T_4 ? _GEN_963 : tag_181; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1734 = _T_4 ? _GEN_964 : tag_182; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1735 = _T_4 ? _GEN_965 : tag_183; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1736 = _T_4 ? _GEN_966 : tag_184; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1737 = _T_4 ? _GEN_967 : tag_185; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1738 = _T_4 ? _GEN_968 : tag_186; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1739 = _T_4 ? _GEN_969 : tag_187; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1740 = _T_4 ? _GEN_970 : tag_188; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1741 = _T_4 ? _GEN_971 : tag_189; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1742 = _T_4 ? _GEN_972 : tag_190; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1743 = _T_4 ? _GEN_973 : tag_191; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1744 = _T_4 ? _GEN_974 : tag_192; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1745 = _T_4 ? _GEN_975 : tag_193; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1746 = _T_4 ? _GEN_976 : tag_194; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1747 = _T_4 ? _GEN_977 : tag_195; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1748 = _T_4 ? _GEN_978 : tag_196; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1749 = _T_4 ? _GEN_979 : tag_197; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1750 = _T_4 ? _GEN_980 : tag_198; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1751 = _T_4 ? _GEN_981 : tag_199; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1752 = _T_4 ? _GEN_982 : tag_200; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1753 = _T_4 ? _GEN_983 : tag_201; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1754 = _T_4 ? _GEN_984 : tag_202; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1755 = _T_4 ? _GEN_985 : tag_203; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1756 = _T_4 ? _GEN_986 : tag_204; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1757 = _T_4 ? _GEN_987 : tag_205; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1758 = _T_4 ? _GEN_988 : tag_206; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1759 = _T_4 ? _GEN_989 : tag_207; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1760 = _T_4 ? _GEN_990 : tag_208; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1761 = _T_4 ? _GEN_991 : tag_209; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1762 = _T_4 ? _GEN_992 : tag_210; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1763 = _T_4 ? _GEN_993 : tag_211; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1764 = _T_4 ? _GEN_994 : tag_212; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1765 = _T_4 ? _GEN_995 : tag_213; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1766 = _T_4 ? _GEN_996 : tag_214; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1767 = _T_4 ? _GEN_997 : tag_215; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1768 = _T_4 ? _GEN_998 : tag_216; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1769 = _T_4 ? _GEN_999 : tag_217; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1770 = _T_4 ? _GEN_1000 : tag_218; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1771 = _T_4 ? _GEN_1001 : tag_219; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1772 = _T_4 ? _GEN_1002 : tag_220; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1773 = _T_4 ? _GEN_1003 : tag_221; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1774 = _T_4 ? _GEN_1004 : tag_222; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1775 = _T_4 ? _GEN_1005 : tag_223; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1776 = _T_4 ? _GEN_1006 : tag_224; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1777 = _T_4 ? _GEN_1007 : tag_225; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1778 = _T_4 ? _GEN_1008 : tag_226; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1779 = _T_4 ? _GEN_1009 : tag_227; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1780 = _T_4 ? _GEN_1010 : tag_228; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1781 = _T_4 ? _GEN_1011 : tag_229; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1782 = _T_4 ? _GEN_1012 : tag_230; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1783 = _T_4 ? _GEN_1013 : tag_231; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1784 = _T_4 ? _GEN_1014 : tag_232; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1785 = _T_4 ? _GEN_1015 : tag_233; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1786 = _T_4 ? _GEN_1016 : tag_234; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1787 = _T_4 ? _GEN_1017 : tag_235; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1788 = _T_4 ? _GEN_1018 : tag_236; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1789 = _T_4 ? _GEN_1019 : tag_237; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1790 = _T_4 ? _GEN_1020 : tag_238; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1791 = _T_4 ? _GEN_1021 : tag_239; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1792 = _T_4 ? _GEN_1022 : tag_240; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1793 = _T_4 ? _GEN_1023 : tag_241; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1794 = _T_4 ? _GEN_1024 : tag_242; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1795 = _T_4 ? _GEN_1025 : tag_243; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1796 = _T_4 ? _GEN_1026 : tag_244; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1797 = _T_4 ? _GEN_1027 : tag_245; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1798 = _T_4 ? _GEN_1028 : tag_246; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1799 = _T_4 ? _GEN_1029 : tag_247; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1800 = _T_4 ? _GEN_1030 : tag_248; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1801 = _T_4 ? _GEN_1031 : tag_249; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1802 = _T_4 ? _GEN_1032 : tag_250; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1803 = _T_4 ? _GEN_1033 : tag_251; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1804 = _T_4 ? _GEN_1034 : tag_252; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1805 = _T_4 ? _GEN_1035 : tag_253; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1806 = _T_4 ? _GEN_1036 : tag_254; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [19:0] _GEN_1807 = _T_4 ? _GEN_1037 : tag_255; // @[Conditional.scala 39:67 Icache.scala 16:24]
  wire [1:0] _GEN_2064 = _T_4 ? 2'h1 : state; // @[Conditional.scala 39:67 Icache.scala 103:25 Icache.scala 25:22]
  wire [31:0] _GEN_2068 = _T_2 ? _GEN_520 : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_2843 = _T_1 ? 1'h0 : _T_2 & _GEN_525; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2845 = _T_1 ? 32'h0 : _GEN_2068; // @[Conditional.scala 39:67]
  S011HD1P_X32Y2D128 req ( // @[Icache.scala 114:19]
    .Q(req_Q),
    .CLK(req_CLK),
    .CEN(req_CEN),
    .WEN(req_WEN),
    .A(req_A),
    .D(req_D)
  );
  assign io_imem_inst_ready = _valid_addr_T & cache_hit; // @[Icache.scala 49:35]
  assign io_imem_inst_read = 2'h3 == req_offset[3:2] ? cache_data_out[127:96] : _inst_read_T_8; // @[Mux.scala 80:57]
  assign io_out_inst_valid = _T ? 1'h0 : _GEN_2843; // @[Conditional.scala 40:58]
  assign io_out_inst_addr = _T ? 32'h0 : _GEN_2845; // @[Conditional.scala 40:58]
  assign req_CLK = clock; // @[Icache.scala 115:14]
  assign req_CEN = 1'h1; // @[Icache.scala 116:14]
  assign req_WEN = cache_wen; // @[Icache.scala 117:14]
  assign req_A = valid_addr[11:4]; // @[Icache.scala 31:28]
  assign req_D = cache_wdata; // @[Icache.scala 119:14]
  always @(posedge clock) begin
    if (reset) begin // @[Icache.scala 16:24]
      tag_0 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_0 <= _GEN_1552;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_1 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_1 <= _GEN_1553;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_2 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_2 <= _GEN_1554;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_3 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_3 <= _GEN_1555;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_4 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_4 <= _GEN_1556;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_5 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_5 <= _GEN_1557;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_6 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_6 <= _GEN_1558;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_7 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_7 <= _GEN_1559;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_8 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_8 <= _GEN_1560;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_9 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_9 <= _GEN_1561;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_10 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_10 <= _GEN_1562;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_11 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_11 <= _GEN_1563;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_12 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_12 <= _GEN_1564;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_13 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_13 <= _GEN_1565;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_14 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_14 <= _GEN_1566;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_15 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_15 <= _GEN_1567;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_16 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_16 <= _GEN_1568;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_17 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_17 <= _GEN_1569;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_18 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_18 <= _GEN_1570;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_19 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_19 <= _GEN_1571;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_20 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_20 <= _GEN_1572;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_21 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_21 <= _GEN_1573;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_22 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_22 <= _GEN_1574;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_23 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_23 <= _GEN_1575;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_24 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_24 <= _GEN_1576;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_25 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_25 <= _GEN_1577;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_26 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_26 <= _GEN_1578;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_27 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_27 <= _GEN_1579;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_28 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_28 <= _GEN_1580;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_29 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_29 <= _GEN_1581;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_30 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_30 <= _GEN_1582;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_31 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_31 <= _GEN_1583;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_32 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_32 <= _GEN_1584;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_33 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_33 <= _GEN_1585;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_34 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_34 <= _GEN_1586;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_35 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_35 <= _GEN_1587;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_36 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_36 <= _GEN_1588;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_37 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_37 <= _GEN_1589;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_38 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_38 <= _GEN_1590;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_39 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_39 <= _GEN_1591;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_40 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_40 <= _GEN_1592;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_41 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_41 <= _GEN_1593;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_42 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_42 <= _GEN_1594;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_43 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_43 <= _GEN_1595;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_44 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_44 <= _GEN_1596;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_45 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_45 <= _GEN_1597;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_46 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_46 <= _GEN_1598;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_47 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_47 <= _GEN_1599;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_48 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_48 <= _GEN_1600;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_49 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_49 <= _GEN_1601;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_50 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_50 <= _GEN_1602;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_51 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_51 <= _GEN_1603;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_52 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_52 <= _GEN_1604;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_53 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_53 <= _GEN_1605;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_54 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_54 <= _GEN_1606;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_55 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_55 <= _GEN_1607;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_56 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_56 <= _GEN_1608;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_57 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_57 <= _GEN_1609;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_58 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_58 <= _GEN_1610;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_59 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_59 <= _GEN_1611;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_60 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_60 <= _GEN_1612;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_61 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_61 <= _GEN_1613;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_62 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_62 <= _GEN_1614;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_63 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_63 <= _GEN_1615;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_64 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_64 <= _GEN_1616;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_65 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_65 <= _GEN_1617;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_66 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_66 <= _GEN_1618;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_67 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_67 <= _GEN_1619;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_68 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_68 <= _GEN_1620;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_69 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_69 <= _GEN_1621;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_70 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_70 <= _GEN_1622;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_71 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_71 <= _GEN_1623;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_72 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_72 <= _GEN_1624;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_73 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_73 <= _GEN_1625;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_74 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_74 <= _GEN_1626;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_75 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_75 <= _GEN_1627;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_76 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_76 <= _GEN_1628;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_77 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_77 <= _GEN_1629;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_78 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_78 <= _GEN_1630;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_79 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_79 <= _GEN_1631;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_80 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_80 <= _GEN_1632;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_81 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_81 <= _GEN_1633;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_82 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_82 <= _GEN_1634;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_83 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_83 <= _GEN_1635;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_84 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_84 <= _GEN_1636;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_85 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_85 <= _GEN_1637;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_86 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_86 <= _GEN_1638;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_87 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_87 <= _GEN_1639;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_88 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_88 <= _GEN_1640;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_89 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_89 <= _GEN_1641;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_90 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_90 <= _GEN_1642;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_91 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_91 <= _GEN_1643;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_92 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_92 <= _GEN_1644;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_93 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_93 <= _GEN_1645;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_94 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_94 <= _GEN_1646;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_95 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_95 <= _GEN_1647;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_96 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_96 <= _GEN_1648;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_97 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_97 <= _GEN_1649;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_98 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_98 <= _GEN_1650;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_99 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_99 <= _GEN_1651;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_100 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_100 <= _GEN_1652;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_101 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_101 <= _GEN_1653;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_102 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_102 <= _GEN_1654;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_103 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_103 <= _GEN_1655;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_104 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_104 <= _GEN_1656;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_105 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_105 <= _GEN_1657;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_106 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_106 <= _GEN_1658;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_107 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_107 <= _GEN_1659;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_108 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_108 <= _GEN_1660;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_109 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_109 <= _GEN_1661;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_110 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_110 <= _GEN_1662;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_111 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_111 <= _GEN_1663;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_112 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_112 <= _GEN_1664;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_113 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_113 <= _GEN_1665;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_114 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_114 <= _GEN_1666;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_115 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_115 <= _GEN_1667;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_116 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_116 <= _GEN_1668;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_117 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_117 <= _GEN_1669;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_118 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_118 <= _GEN_1670;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_119 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_119 <= _GEN_1671;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_120 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_120 <= _GEN_1672;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_121 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_121 <= _GEN_1673;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_122 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_122 <= _GEN_1674;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_123 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_123 <= _GEN_1675;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_124 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_124 <= _GEN_1676;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_125 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_125 <= _GEN_1677;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_126 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_126 <= _GEN_1678;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_127 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_127 <= _GEN_1679;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_128 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_128 <= _GEN_1680;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_129 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_129 <= _GEN_1681;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_130 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_130 <= _GEN_1682;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_131 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_131 <= _GEN_1683;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_132 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_132 <= _GEN_1684;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_133 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_133 <= _GEN_1685;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_134 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_134 <= _GEN_1686;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_135 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_135 <= _GEN_1687;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_136 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_136 <= _GEN_1688;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_137 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_137 <= _GEN_1689;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_138 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_138 <= _GEN_1690;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_139 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_139 <= _GEN_1691;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_140 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_140 <= _GEN_1692;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_141 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_141 <= _GEN_1693;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_142 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_142 <= _GEN_1694;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_143 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_143 <= _GEN_1695;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_144 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_144 <= _GEN_1696;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_145 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_145 <= _GEN_1697;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_146 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_146 <= _GEN_1698;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_147 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_147 <= _GEN_1699;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_148 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_148 <= _GEN_1700;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_149 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_149 <= _GEN_1701;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_150 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_150 <= _GEN_1702;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_151 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_151 <= _GEN_1703;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_152 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_152 <= _GEN_1704;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_153 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_153 <= _GEN_1705;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_154 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_154 <= _GEN_1706;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_155 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_155 <= _GEN_1707;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_156 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_156 <= _GEN_1708;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_157 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_157 <= _GEN_1709;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_158 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_158 <= _GEN_1710;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_159 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_159 <= _GEN_1711;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_160 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_160 <= _GEN_1712;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_161 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_161 <= _GEN_1713;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_162 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_162 <= _GEN_1714;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_163 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_163 <= _GEN_1715;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_164 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_164 <= _GEN_1716;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_165 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_165 <= _GEN_1717;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_166 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_166 <= _GEN_1718;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_167 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_167 <= _GEN_1719;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_168 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_168 <= _GEN_1720;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_169 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_169 <= _GEN_1721;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_170 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_170 <= _GEN_1722;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_171 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_171 <= _GEN_1723;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_172 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_172 <= _GEN_1724;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_173 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_173 <= _GEN_1725;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_174 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_174 <= _GEN_1726;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_175 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_175 <= _GEN_1727;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_176 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_176 <= _GEN_1728;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_177 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_177 <= _GEN_1729;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_178 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_178 <= _GEN_1730;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_179 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_179 <= _GEN_1731;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_180 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_180 <= _GEN_1732;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_181 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_181 <= _GEN_1733;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_182 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_182 <= _GEN_1734;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_183 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_183 <= _GEN_1735;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_184 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_184 <= _GEN_1736;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_185 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_185 <= _GEN_1737;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_186 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_186 <= _GEN_1738;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_187 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_187 <= _GEN_1739;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_188 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_188 <= _GEN_1740;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_189 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_189 <= _GEN_1741;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_190 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_190 <= _GEN_1742;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_191 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_191 <= _GEN_1743;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_192 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_192 <= _GEN_1744;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_193 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_193 <= _GEN_1745;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_194 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_194 <= _GEN_1746;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_195 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_195 <= _GEN_1747;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_196 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_196 <= _GEN_1748;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_197 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_197 <= _GEN_1749;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_198 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_198 <= _GEN_1750;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_199 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_199 <= _GEN_1751;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_200 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_200 <= _GEN_1752;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_201 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_201 <= _GEN_1753;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_202 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_202 <= _GEN_1754;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_203 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_203 <= _GEN_1755;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_204 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_204 <= _GEN_1756;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_205 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_205 <= _GEN_1757;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_206 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_206 <= _GEN_1758;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_207 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_207 <= _GEN_1759;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_208 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_208 <= _GEN_1760;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_209 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_209 <= _GEN_1761;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_210 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_210 <= _GEN_1762;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_211 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_211 <= _GEN_1763;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_212 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_212 <= _GEN_1764;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_213 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_213 <= _GEN_1765;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_214 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_214 <= _GEN_1766;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_215 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_215 <= _GEN_1767;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_216 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_216 <= _GEN_1768;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_217 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_217 <= _GEN_1769;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_218 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_218 <= _GEN_1770;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_219 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_219 <= _GEN_1771;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_220 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_220 <= _GEN_1772;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_221 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_221 <= _GEN_1773;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_222 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_222 <= _GEN_1774;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_223 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_223 <= _GEN_1775;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_224 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_224 <= _GEN_1776;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_225 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_225 <= _GEN_1777;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_226 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_226 <= _GEN_1778;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_227 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_227 <= _GEN_1779;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_228 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_228 <= _GEN_1780;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_229 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_229 <= _GEN_1781;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_230 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_230 <= _GEN_1782;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_231 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_231 <= _GEN_1783;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_232 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_232 <= _GEN_1784;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_233 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_233 <= _GEN_1785;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_234 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_234 <= _GEN_1786;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_235 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_235 <= _GEN_1787;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_236 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_236 <= _GEN_1788;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_237 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_237 <= _GEN_1789;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_238 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_238 <= _GEN_1790;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_239 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_239 <= _GEN_1791;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_240 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_240 <= _GEN_1792;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_241 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_241 <= _GEN_1793;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_242 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_242 <= _GEN_1794;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_243 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_243 <= _GEN_1795;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_244 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_244 <= _GEN_1796;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_245 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_245 <= _GEN_1797;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_246 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_246 <= _GEN_1798;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_247 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_247 <= _GEN_1799;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_248 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_248 <= _GEN_1800;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_249 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_249 <= _GEN_1801;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_250 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_250 <= _GEN_1802;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_251 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_251 <= _GEN_1803;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_252 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_252 <= _GEN_1804;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_253 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_253 <= _GEN_1805;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_254 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_254 <= _GEN_1806;
        end
      end
    end
    if (reset) begin // @[Icache.scala 16:24]
      tag_255 <= 20'h0; // @[Icache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          tag_255 <= _GEN_1807;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_0 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_0 <= _GEN_1296;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_1 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_1 <= _GEN_1297;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_2 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_2 <= _GEN_1298;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_3 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_3 <= _GEN_1299;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_4 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_4 <= _GEN_1300;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_5 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_5 <= _GEN_1301;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_6 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_6 <= _GEN_1302;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_7 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_7 <= _GEN_1303;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_8 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_8 <= _GEN_1304;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_9 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_9 <= _GEN_1305;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_10 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_10 <= _GEN_1306;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_11 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_11 <= _GEN_1307;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_12 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_12 <= _GEN_1308;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_13 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_13 <= _GEN_1309;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_14 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_14 <= _GEN_1310;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_15 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_15 <= _GEN_1311;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_16 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_16 <= _GEN_1312;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_17 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_17 <= _GEN_1313;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_18 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_18 <= _GEN_1314;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_19 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_19 <= _GEN_1315;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_20 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_20 <= _GEN_1316;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_21 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_21 <= _GEN_1317;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_22 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_22 <= _GEN_1318;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_23 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_23 <= _GEN_1319;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_24 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_24 <= _GEN_1320;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_25 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_25 <= _GEN_1321;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_26 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_26 <= _GEN_1322;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_27 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_27 <= _GEN_1323;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_28 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_28 <= _GEN_1324;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_29 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_29 <= _GEN_1325;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_30 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_30 <= _GEN_1326;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_31 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_31 <= _GEN_1327;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_32 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_32 <= _GEN_1328;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_33 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_33 <= _GEN_1329;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_34 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_34 <= _GEN_1330;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_35 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_35 <= _GEN_1331;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_36 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_36 <= _GEN_1332;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_37 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_37 <= _GEN_1333;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_38 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_38 <= _GEN_1334;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_39 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_39 <= _GEN_1335;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_40 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_40 <= _GEN_1336;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_41 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_41 <= _GEN_1337;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_42 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_42 <= _GEN_1338;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_43 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_43 <= _GEN_1339;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_44 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_44 <= _GEN_1340;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_45 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_45 <= _GEN_1341;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_46 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_46 <= _GEN_1342;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_47 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_47 <= _GEN_1343;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_48 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_48 <= _GEN_1344;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_49 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_49 <= _GEN_1345;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_50 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_50 <= _GEN_1346;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_51 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_51 <= _GEN_1347;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_52 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_52 <= _GEN_1348;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_53 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_53 <= _GEN_1349;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_54 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_54 <= _GEN_1350;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_55 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_55 <= _GEN_1351;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_56 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_56 <= _GEN_1352;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_57 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_57 <= _GEN_1353;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_58 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_58 <= _GEN_1354;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_59 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_59 <= _GEN_1355;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_60 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_60 <= _GEN_1356;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_61 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_61 <= _GEN_1357;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_62 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_62 <= _GEN_1358;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_63 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_63 <= _GEN_1359;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_64 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_64 <= _GEN_1360;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_65 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_65 <= _GEN_1361;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_66 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_66 <= _GEN_1362;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_67 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_67 <= _GEN_1363;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_68 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_68 <= _GEN_1364;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_69 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_69 <= _GEN_1365;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_70 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_70 <= _GEN_1366;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_71 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_71 <= _GEN_1367;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_72 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_72 <= _GEN_1368;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_73 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_73 <= _GEN_1369;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_74 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_74 <= _GEN_1370;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_75 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_75 <= _GEN_1371;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_76 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_76 <= _GEN_1372;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_77 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_77 <= _GEN_1373;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_78 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_78 <= _GEN_1374;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_79 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_79 <= _GEN_1375;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_80 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_80 <= _GEN_1376;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_81 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_81 <= _GEN_1377;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_82 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_82 <= _GEN_1378;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_83 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_83 <= _GEN_1379;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_84 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_84 <= _GEN_1380;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_85 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_85 <= _GEN_1381;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_86 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_86 <= _GEN_1382;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_87 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_87 <= _GEN_1383;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_88 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_88 <= _GEN_1384;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_89 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_89 <= _GEN_1385;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_90 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_90 <= _GEN_1386;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_91 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_91 <= _GEN_1387;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_92 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_92 <= _GEN_1388;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_93 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_93 <= _GEN_1389;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_94 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_94 <= _GEN_1390;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_95 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_95 <= _GEN_1391;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_96 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_96 <= _GEN_1392;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_97 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_97 <= _GEN_1393;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_98 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_98 <= _GEN_1394;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_99 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_99 <= _GEN_1395;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_100 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_100 <= _GEN_1396;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_101 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_101 <= _GEN_1397;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_102 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_102 <= _GEN_1398;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_103 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_103 <= _GEN_1399;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_104 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_104 <= _GEN_1400;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_105 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_105 <= _GEN_1401;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_106 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_106 <= _GEN_1402;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_107 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_107 <= _GEN_1403;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_108 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_108 <= _GEN_1404;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_109 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_109 <= _GEN_1405;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_110 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_110 <= _GEN_1406;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_111 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_111 <= _GEN_1407;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_112 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_112 <= _GEN_1408;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_113 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_113 <= _GEN_1409;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_114 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_114 <= _GEN_1410;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_115 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_115 <= _GEN_1411;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_116 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_116 <= _GEN_1412;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_117 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_117 <= _GEN_1413;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_118 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_118 <= _GEN_1414;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_119 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_119 <= _GEN_1415;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_120 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_120 <= _GEN_1416;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_121 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_121 <= _GEN_1417;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_122 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_122 <= _GEN_1418;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_123 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_123 <= _GEN_1419;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_124 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_124 <= _GEN_1420;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_125 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_125 <= _GEN_1421;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_126 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_126 <= _GEN_1422;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_127 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_127 <= _GEN_1423;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_128 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_128 <= _GEN_1424;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_129 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_129 <= _GEN_1425;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_130 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_130 <= _GEN_1426;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_131 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_131 <= _GEN_1427;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_132 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_132 <= _GEN_1428;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_133 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_133 <= _GEN_1429;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_134 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_134 <= _GEN_1430;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_135 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_135 <= _GEN_1431;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_136 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_136 <= _GEN_1432;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_137 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_137 <= _GEN_1433;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_138 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_138 <= _GEN_1434;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_139 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_139 <= _GEN_1435;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_140 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_140 <= _GEN_1436;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_141 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_141 <= _GEN_1437;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_142 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_142 <= _GEN_1438;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_143 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_143 <= _GEN_1439;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_144 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_144 <= _GEN_1440;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_145 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_145 <= _GEN_1441;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_146 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_146 <= _GEN_1442;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_147 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_147 <= _GEN_1443;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_148 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_148 <= _GEN_1444;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_149 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_149 <= _GEN_1445;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_150 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_150 <= _GEN_1446;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_151 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_151 <= _GEN_1447;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_152 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_152 <= _GEN_1448;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_153 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_153 <= _GEN_1449;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_154 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_154 <= _GEN_1450;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_155 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_155 <= _GEN_1451;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_156 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_156 <= _GEN_1452;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_157 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_157 <= _GEN_1453;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_158 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_158 <= _GEN_1454;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_159 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_159 <= _GEN_1455;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_160 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_160 <= _GEN_1456;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_161 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_161 <= _GEN_1457;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_162 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_162 <= _GEN_1458;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_163 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_163 <= _GEN_1459;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_164 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_164 <= _GEN_1460;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_165 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_165 <= _GEN_1461;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_166 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_166 <= _GEN_1462;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_167 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_167 <= _GEN_1463;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_168 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_168 <= _GEN_1464;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_169 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_169 <= _GEN_1465;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_170 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_170 <= _GEN_1466;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_171 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_171 <= _GEN_1467;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_172 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_172 <= _GEN_1468;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_173 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_173 <= _GEN_1469;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_174 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_174 <= _GEN_1470;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_175 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_175 <= _GEN_1471;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_176 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_176 <= _GEN_1472;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_177 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_177 <= _GEN_1473;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_178 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_178 <= _GEN_1474;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_179 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_179 <= _GEN_1475;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_180 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_180 <= _GEN_1476;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_181 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_181 <= _GEN_1477;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_182 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_182 <= _GEN_1478;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_183 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_183 <= _GEN_1479;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_184 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_184 <= _GEN_1480;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_185 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_185 <= _GEN_1481;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_186 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_186 <= _GEN_1482;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_187 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_187 <= _GEN_1483;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_188 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_188 <= _GEN_1484;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_189 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_189 <= _GEN_1485;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_190 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_190 <= _GEN_1486;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_191 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_191 <= _GEN_1487;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_192 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_192 <= _GEN_1488;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_193 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_193 <= _GEN_1489;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_194 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_194 <= _GEN_1490;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_195 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_195 <= _GEN_1491;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_196 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_196 <= _GEN_1492;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_197 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_197 <= _GEN_1493;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_198 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_198 <= _GEN_1494;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_199 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_199 <= _GEN_1495;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_200 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_200 <= _GEN_1496;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_201 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_201 <= _GEN_1497;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_202 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_202 <= _GEN_1498;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_203 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_203 <= _GEN_1499;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_204 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_204 <= _GEN_1500;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_205 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_205 <= _GEN_1501;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_206 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_206 <= _GEN_1502;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_207 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_207 <= _GEN_1503;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_208 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_208 <= _GEN_1504;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_209 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_209 <= _GEN_1505;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_210 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_210 <= _GEN_1506;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_211 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_211 <= _GEN_1507;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_212 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_212 <= _GEN_1508;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_213 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_213 <= _GEN_1509;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_214 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_214 <= _GEN_1510;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_215 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_215 <= _GEN_1511;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_216 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_216 <= _GEN_1512;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_217 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_217 <= _GEN_1513;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_218 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_218 <= _GEN_1514;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_219 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_219 <= _GEN_1515;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_220 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_220 <= _GEN_1516;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_221 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_221 <= _GEN_1517;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_222 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_222 <= _GEN_1518;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_223 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_223 <= _GEN_1519;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_224 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_224 <= _GEN_1520;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_225 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_225 <= _GEN_1521;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_226 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_226 <= _GEN_1522;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_227 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_227 <= _GEN_1523;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_228 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_228 <= _GEN_1524;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_229 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_229 <= _GEN_1525;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_230 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_230 <= _GEN_1526;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_231 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_231 <= _GEN_1527;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_232 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_232 <= _GEN_1528;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_233 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_233 <= _GEN_1529;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_234 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_234 <= _GEN_1530;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_235 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_235 <= _GEN_1531;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_236 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_236 <= _GEN_1532;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_237 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_237 <= _GEN_1533;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_238 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_238 <= _GEN_1534;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_239 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_239 <= _GEN_1535;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_240 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_240 <= _GEN_1536;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_241 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_241 <= _GEN_1537;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_242 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_242 <= _GEN_1538;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_243 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_243 <= _GEN_1539;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_244 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_244 <= _GEN_1540;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_245 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_245 <= _GEN_1541;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_246 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_246 <= _GEN_1542;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_247 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_247 <= _GEN_1543;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_248 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_248 <= _GEN_1544;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_249 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_249 <= _GEN_1545;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_250 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_250 <= _GEN_1546;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_251 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_251 <= _GEN_1547;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_252 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_252 <= _GEN_1548;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_253 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_253 <= _GEN_1549;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_254 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_254 <= _GEN_1550;
        end
      end
    end
    if (reset) begin // @[Icache.scala 17:24]
      valid_255 <= 1'h0; // @[Icache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_2)) begin // @[Conditional.scala 39:67]
          valid_255 <= _GEN_1551;
        end
      end
    end
    if (reset) begin // @[Icache.scala 25:22]
      state <= 2'h0; // @[Icache.scala 25:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_imem_inst_valid) begin // @[Icache.scala 57:28]
        state <= 2'h1; // @[Icache.scala 58:15]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (io_imem_inst_valid) begin // @[Icache.scala 63:28]
        state <= _GEN_514;
      end else begin
        state <= 2'h0; // @[Icache.scala 74:15]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      state <= _GEN_517;
    end else begin
      state <= _GEN_2064;
    end
    if (reset) begin // @[Icache.scala 27:27]
      req_addr <= 32'h0; // @[Icache.scala 27:27]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (io_imem_inst_valid) begin // @[Icache.scala 63:28]
          req_addr <= io_imem_inst_addr;
        end
      end
    end
    if (reset) begin // @[Icache.scala 51:28]
      cache_fill <= 1'h0; // @[Icache.scala 51:28]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          cache_fill <= _GEN_522;
        end else begin
          cache_fill <= _GEN_1294;
        end
      end
    end
    if (reset) begin // @[Icache.scala 52:28]
      cache_wen <= 1'h0; // @[Icache.scala 52:28]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          cache_wen <= _GEN_523;
        end else begin
          cache_wen <= _GEN_1295;
        end
      end
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_wdata <= 128'h0; // @[Icache.scala 53:28]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[Conditional.scala 39:67]
          cache_wdata <= _GEN_524;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_0 = _RAND_0[19:0];
  _RAND_1 = {1{`RANDOM}};
  tag_1 = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  tag_2 = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  tag_3 = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  tag_4 = _RAND_4[19:0];
  _RAND_5 = {1{`RANDOM}};
  tag_5 = _RAND_5[19:0];
  _RAND_6 = {1{`RANDOM}};
  tag_6 = _RAND_6[19:0];
  _RAND_7 = {1{`RANDOM}};
  tag_7 = _RAND_7[19:0];
  _RAND_8 = {1{`RANDOM}};
  tag_8 = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  tag_9 = _RAND_9[19:0];
  _RAND_10 = {1{`RANDOM}};
  tag_10 = _RAND_10[19:0];
  _RAND_11 = {1{`RANDOM}};
  tag_11 = _RAND_11[19:0];
  _RAND_12 = {1{`RANDOM}};
  tag_12 = _RAND_12[19:0];
  _RAND_13 = {1{`RANDOM}};
  tag_13 = _RAND_13[19:0];
  _RAND_14 = {1{`RANDOM}};
  tag_14 = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  tag_15 = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  tag_16 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  tag_17 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  tag_18 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  tag_19 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  tag_20 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  tag_21 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  tag_22 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  tag_23 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  tag_24 = _RAND_24[19:0];
  _RAND_25 = {1{`RANDOM}};
  tag_25 = _RAND_25[19:0];
  _RAND_26 = {1{`RANDOM}};
  tag_26 = _RAND_26[19:0];
  _RAND_27 = {1{`RANDOM}};
  tag_27 = _RAND_27[19:0];
  _RAND_28 = {1{`RANDOM}};
  tag_28 = _RAND_28[19:0];
  _RAND_29 = {1{`RANDOM}};
  tag_29 = _RAND_29[19:0];
  _RAND_30 = {1{`RANDOM}};
  tag_30 = _RAND_30[19:0];
  _RAND_31 = {1{`RANDOM}};
  tag_31 = _RAND_31[19:0];
  _RAND_32 = {1{`RANDOM}};
  tag_32 = _RAND_32[19:0];
  _RAND_33 = {1{`RANDOM}};
  tag_33 = _RAND_33[19:0];
  _RAND_34 = {1{`RANDOM}};
  tag_34 = _RAND_34[19:0];
  _RAND_35 = {1{`RANDOM}};
  tag_35 = _RAND_35[19:0];
  _RAND_36 = {1{`RANDOM}};
  tag_36 = _RAND_36[19:0];
  _RAND_37 = {1{`RANDOM}};
  tag_37 = _RAND_37[19:0];
  _RAND_38 = {1{`RANDOM}};
  tag_38 = _RAND_38[19:0];
  _RAND_39 = {1{`RANDOM}};
  tag_39 = _RAND_39[19:0];
  _RAND_40 = {1{`RANDOM}};
  tag_40 = _RAND_40[19:0];
  _RAND_41 = {1{`RANDOM}};
  tag_41 = _RAND_41[19:0];
  _RAND_42 = {1{`RANDOM}};
  tag_42 = _RAND_42[19:0];
  _RAND_43 = {1{`RANDOM}};
  tag_43 = _RAND_43[19:0];
  _RAND_44 = {1{`RANDOM}};
  tag_44 = _RAND_44[19:0];
  _RAND_45 = {1{`RANDOM}};
  tag_45 = _RAND_45[19:0];
  _RAND_46 = {1{`RANDOM}};
  tag_46 = _RAND_46[19:0];
  _RAND_47 = {1{`RANDOM}};
  tag_47 = _RAND_47[19:0];
  _RAND_48 = {1{`RANDOM}};
  tag_48 = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  tag_49 = _RAND_49[19:0];
  _RAND_50 = {1{`RANDOM}};
  tag_50 = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  tag_51 = _RAND_51[19:0];
  _RAND_52 = {1{`RANDOM}};
  tag_52 = _RAND_52[19:0];
  _RAND_53 = {1{`RANDOM}};
  tag_53 = _RAND_53[19:0];
  _RAND_54 = {1{`RANDOM}};
  tag_54 = _RAND_54[19:0];
  _RAND_55 = {1{`RANDOM}};
  tag_55 = _RAND_55[19:0];
  _RAND_56 = {1{`RANDOM}};
  tag_56 = _RAND_56[19:0];
  _RAND_57 = {1{`RANDOM}};
  tag_57 = _RAND_57[19:0];
  _RAND_58 = {1{`RANDOM}};
  tag_58 = _RAND_58[19:0];
  _RAND_59 = {1{`RANDOM}};
  tag_59 = _RAND_59[19:0];
  _RAND_60 = {1{`RANDOM}};
  tag_60 = _RAND_60[19:0];
  _RAND_61 = {1{`RANDOM}};
  tag_61 = _RAND_61[19:0];
  _RAND_62 = {1{`RANDOM}};
  tag_62 = _RAND_62[19:0];
  _RAND_63 = {1{`RANDOM}};
  tag_63 = _RAND_63[19:0];
  _RAND_64 = {1{`RANDOM}};
  tag_64 = _RAND_64[19:0];
  _RAND_65 = {1{`RANDOM}};
  tag_65 = _RAND_65[19:0];
  _RAND_66 = {1{`RANDOM}};
  tag_66 = _RAND_66[19:0];
  _RAND_67 = {1{`RANDOM}};
  tag_67 = _RAND_67[19:0];
  _RAND_68 = {1{`RANDOM}};
  tag_68 = _RAND_68[19:0];
  _RAND_69 = {1{`RANDOM}};
  tag_69 = _RAND_69[19:0];
  _RAND_70 = {1{`RANDOM}};
  tag_70 = _RAND_70[19:0];
  _RAND_71 = {1{`RANDOM}};
  tag_71 = _RAND_71[19:0];
  _RAND_72 = {1{`RANDOM}};
  tag_72 = _RAND_72[19:0];
  _RAND_73 = {1{`RANDOM}};
  tag_73 = _RAND_73[19:0];
  _RAND_74 = {1{`RANDOM}};
  tag_74 = _RAND_74[19:0];
  _RAND_75 = {1{`RANDOM}};
  tag_75 = _RAND_75[19:0];
  _RAND_76 = {1{`RANDOM}};
  tag_76 = _RAND_76[19:0];
  _RAND_77 = {1{`RANDOM}};
  tag_77 = _RAND_77[19:0];
  _RAND_78 = {1{`RANDOM}};
  tag_78 = _RAND_78[19:0];
  _RAND_79 = {1{`RANDOM}};
  tag_79 = _RAND_79[19:0];
  _RAND_80 = {1{`RANDOM}};
  tag_80 = _RAND_80[19:0];
  _RAND_81 = {1{`RANDOM}};
  tag_81 = _RAND_81[19:0];
  _RAND_82 = {1{`RANDOM}};
  tag_82 = _RAND_82[19:0];
  _RAND_83 = {1{`RANDOM}};
  tag_83 = _RAND_83[19:0];
  _RAND_84 = {1{`RANDOM}};
  tag_84 = _RAND_84[19:0];
  _RAND_85 = {1{`RANDOM}};
  tag_85 = _RAND_85[19:0];
  _RAND_86 = {1{`RANDOM}};
  tag_86 = _RAND_86[19:0];
  _RAND_87 = {1{`RANDOM}};
  tag_87 = _RAND_87[19:0];
  _RAND_88 = {1{`RANDOM}};
  tag_88 = _RAND_88[19:0];
  _RAND_89 = {1{`RANDOM}};
  tag_89 = _RAND_89[19:0];
  _RAND_90 = {1{`RANDOM}};
  tag_90 = _RAND_90[19:0];
  _RAND_91 = {1{`RANDOM}};
  tag_91 = _RAND_91[19:0];
  _RAND_92 = {1{`RANDOM}};
  tag_92 = _RAND_92[19:0];
  _RAND_93 = {1{`RANDOM}};
  tag_93 = _RAND_93[19:0];
  _RAND_94 = {1{`RANDOM}};
  tag_94 = _RAND_94[19:0];
  _RAND_95 = {1{`RANDOM}};
  tag_95 = _RAND_95[19:0];
  _RAND_96 = {1{`RANDOM}};
  tag_96 = _RAND_96[19:0];
  _RAND_97 = {1{`RANDOM}};
  tag_97 = _RAND_97[19:0];
  _RAND_98 = {1{`RANDOM}};
  tag_98 = _RAND_98[19:0];
  _RAND_99 = {1{`RANDOM}};
  tag_99 = _RAND_99[19:0];
  _RAND_100 = {1{`RANDOM}};
  tag_100 = _RAND_100[19:0];
  _RAND_101 = {1{`RANDOM}};
  tag_101 = _RAND_101[19:0];
  _RAND_102 = {1{`RANDOM}};
  tag_102 = _RAND_102[19:0];
  _RAND_103 = {1{`RANDOM}};
  tag_103 = _RAND_103[19:0];
  _RAND_104 = {1{`RANDOM}};
  tag_104 = _RAND_104[19:0];
  _RAND_105 = {1{`RANDOM}};
  tag_105 = _RAND_105[19:0];
  _RAND_106 = {1{`RANDOM}};
  tag_106 = _RAND_106[19:0];
  _RAND_107 = {1{`RANDOM}};
  tag_107 = _RAND_107[19:0];
  _RAND_108 = {1{`RANDOM}};
  tag_108 = _RAND_108[19:0];
  _RAND_109 = {1{`RANDOM}};
  tag_109 = _RAND_109[19:0];
  _RAND_110 = {1{`RANDOM}};
  tag_110 = _RAND_110[19:0];
  _RAND_111 = {1{`RANDOM}};
  tag_111 = _RAND_111[19:0];
  _RAND_112 = {1{`RANDOM}};
  tag_112 = _RAND_112[19:0];
  _RAND_113 = {1{`RANDOM}};
  tag_113 = _RAND_113[19:0];
  _RAND_114 = {1{`RANDOM}};
  tag_114 = _RAND_114[19:0];
  _RAND_115 = {1{`RANDOM}};
  tag_115 = _RAND_115[19:0];
  _RAND_116 = {1{`RANDOM}};
  tag_116 = _RAND_116[19:0];
  _RAND_117 = {1{`RANDOM}};
  tag_117 = _RAND_117[19:0];
  _RAND_118 = {1{`RANDOM}};
  tag_118 = _RAND_118[19:0];
  _RAND_119 = {1{`RANDOM}};
  tag_119 = _RAND_119[19:0];
  _RAND_120 = {1{`RANDOM}};
  tag_120 = _RAND_120[19:0];
  _RAND_121 = {1{`RANDOM}};
  tag_121 = _RAND_121[19:0];
  _RAND_122 = {1{`RANDOM}};
  tag_122 = _RAND_122[19:0];
  _RAND_123 = {1{`RANDOM}};
  tag_123 = _RAND_123[19:0];
  _RAND_124 = {1{`RANDOM}};
  tag_124 = _RAND_124[19:0];
  _RAND_125 = {1{`RANDOM}};
  tag_125 = _RAND_125[19:0];
  _RAND_126 = {1{`RANDOM}};
  tag_126 = _RAND_126[19:0];
  _RAND_127 = {1{`RANDOM}};
  tag_127 = _RAND_127[19:0];
  _RAND_128 = {1{`RANDOM}};
  tag_128 = _RAND_128[19:0];
  _RAND_129 = {1{`RANDOM}};
  tag_129 = _RAND_129[19:0];
  _RAND_130 = {1{`RANDOM}};
  tag_130 = _RAND_130[19:0];
  _RAND_131 = {1{`RANDOM}};
  tag_131 = _RAND_131[19:0];
  _RAND_132 = {1{`RANDOM}};
  tag_132 = _RAND_132[19:0];
  _RAND_133 = {1{`RANDOM}};
  tag_133 = _RAND_133[19:0];
  _RAND_134 = {1{`RANDOM}};
  tag_134 = _RAND_134[19:0];
  _RAND_135 = {1{`RANDOM}};
  tag_135 = _RAND_135[19:0];
  _RAND_136 = {1{`RANDOM}};
  tag_136 = _RAND_136[19:0];
  _RAND_137 = {1{`RANDOM}};
  tag_137 = _RAND_137[19:0];
  _RAND_138 = {1{`RANDOM}};
  tag_138 = _RAND_138[19:0];
  _RAND_139 = {1{`RANDOM}};
  tag_139 = _RAND_139[19:0];
  _RAND_140 = {1{`RANDOM}};
  tag_140 = _RAND_140[19:0];
  _RAND_141 = {1{`RANDOM}};
  tag_141 = _RAND_141[19:0];
  _RAND_142 = {1{`RANDOM}};
  tag_142 = _RAND_142[19:0];
  _RAND_143 = {1{`RANDOM}};
  tag_143 = _RAND_143[19:0];
  _RAND_144 = {1{`RANDOM}};
  tag_144 = _RAND_144[19:0];
  _RAND_145 = {1{`RANDOM}};
  tag_145 = _RAND_145[19:0];
  _RAND_146 = {1{`RANDOM}};
  tag_146 = _RAND_146[19:0];
  _RAND_147 = {1{`RANDOM}};
  tag_147 = _RAND_147[19:0];
  _RAND_148 = {1{`RANDOM}};
  tag_148 = _RAND_148[19:0];
  _RAND_149 = {1{`RANDOM}};
  tag_149 = _RAND_149[19:0];
  _RAND_150 = {1{`RANDOM}};
  tag_150 = _RAND_150[19:0];
  _RAND_151 = {1{`RANDOM}};
  tag_151 = _RAND_151[19:0];
  _RAND_152 = {1{`RANDOM}};
  tag_152 = _RAND_152[19:0];
  _RAND_153 = {1{`RANDOM}};
  tag_153 = _RAND_153[19:0];
  _RAND_154 = {1{`RANDOM}};
  tag_154 = _RAND_154[19:0];
  _RAND_155 = {1{`RANDOM}};
  tag_155 = _RAND_155[19:0];
  _RAND_156 = {1{`RANDOM}};
  tag_156 = _RAND_156[19:0];
  _RAND_157 = {1{`RANDOM}};
  tag_157 = _RAND_157[19:0];
  _RAND_158 = {1{`RANDOM}};
  tag_158 = _RAND_158[19:0];
  _RAND_159 = {1{`RANDOM}};
  tag_159 = _RAND_159[19:0];
  _RAND_160 = {1{`RANDOM}};
  tag_160 = _RAND_160[19:0];
  _RAND_161 = {1{`RANDOM}};
  tag_161 = _RAND_161[19:0];
  _RAND_162 = {1{`RANDOM}};
  tag_162 = _RAND_162[19:0];
  _RAND_163 = {1{`RANDOM}};
  tag_163 = _RAND_163[19:0];
  _RAND_164 = {1{`RANDOM}};
  tag_164 = _RAND_164[19:0];
  _RAND_165 = {1{`RANDOM}};
  tag_165 = _RAND_165[19:0];
  _RAND_166 = {1{`RANDOM}};
  tag_166 = _RAND_166[19:0];
  _RAND_167 = {1{`RANDOM}};
  tag_167 = _RAND_167[19:0];
  _RAND_168 = {1{`RANDOM}};
  tag_168 = _RAND_168[19:0];
  _RAND_169 = {1{`RANDOM}};
  tag_169 = _RAND_169[19:0];
  _RAND_170 = {1{`RANDOM}};
  tag_170 = _RAND_170[19:0];
  _RAND_171 = {1{`RANDOM}};
  tag_171 = _RAND_171[19:0];
  _RAND_172 = {1{`RANDOM}};
  tag_172 = _RAND_172[19:0];
  _RAND_173 = {1{`RANDOM}};
  tag_173 = _RAND_173[19:0];
  _RAND_174 = {1{`RANDOM}};
  tag_174 = _RAND_174[19:0];
  _RAND_175 = {1{`RANDOM}};
  tag_175 = _RAND_175[19:0];
  _RAND_176 = {1{`RANDOM}};
  tag_176 = _RAND_176[19:0];
  _RAND_177 = {1{`RANDOM}};
  tag_177 = _RAND_177[19:0];
  _RAND_178 = {1{`RANDOM}};
  tag_178 = _RAND_178[19:0];
  _RAND_179 = {1{`RANDOM}};
  tag_179 = _RAND_179[19:0];
  _RAND_180 = {1{`RANDOM}};
  tag_180 = _RAND_180[19:0];
  _RAND_181 = {1{`RANDOM}};
  tag_181 = _RAND_181[19:0];
  _RAND_182 = {1{`RANDOM}};
  tag_182 = _RAND_182[19:0];
  _RAND_183 = {1{`RANDOM}};
  tag_183 = _RAND_183[19:0];
  _RAND_184 = {1{`RANDOM}};
  tag_184 = _RAND_184[19:0];
  _RAND_185 = {1{`RANDOM}};
  tag_185 = _RAND_185[19:0];
  _RAND_186 = {1{`RANDOM}};
  tag_186 = _RAND_186[19:0];
  _RAND_187 = {1{`RANDOM}};
  tag_187 = _RAND_187[19:0];
  _RAND_188 = {1{`RANDOM}};
  tag_188 = _RAND_188[19:0];
  _RAND_189 = {1{`RANDOM}};
  tag_189 = _RAND_189[19:0];
  _RAND_190 = {1{`RANDOM}};
  tag_190 = _RAND_190[19:0];
  _RAND_191 = {1{`RANDOM}};
  tag_191 = _RAND_191[19:0];
  _RAND_192 = {1{`RANDOM}};
  tag_192 = _RAND_192[19:0];
  _RAND_193 = {1{`RANDOM}};
  tag_193 = _RAND_193[19:0];
  _RAND_194 = {1{`RANDOM}};
  tag_194 = _RAND_194[19:0];
  _RAND_195 = {1{`RANDOM}};
  tag_195 = _RAND_195[19:0];
  _RAND_196 = {1{`RANDOM}};
  tag_196 = _RAND_196[19:0];
  _RAND_197 = {1{`RANDOM}};
  tag_197 = _RAND_197[19:0];
  _RAND_198 = {1{`RANDOM}};
  tag_198 = _RAND_198[19:0];
  _RAND_199 = {1{`RANDOM}};
  tag_199 = _RAND_199[19:0];
  _RAND_200 = {1{`RANDOM}};
  tag_200 = _RAND_200[19:0];
  _RAND_201 = {1{`RANDOM}};
  tag_201 = _RAND_201[19:0];
  _RAND_202 = {1{`RANDOM}};
  tag_202 = _RAND_202[19:0];
  _RAND_203 = {1{`RANDOM}};
  tag_203 = _RAND_203[19:0];
  _RAND_204 = {1{`RANDOM}};
  tag_204 = _RAND_204[19:0];
  _RAND_205 = {1{`RANDOM}};
  tag_205 = _RAND_205[19:0];
  _RAND_206 = {1{`RANDOM}};
  tag_206 = _RAND_206[19:0];
  _RAND_207 = {1{`RANDOM}};
  tag_207 = _RAND_207[19:0];
  _RAND_208 = {1{`RANDOM}};
  tag_208 = _RAND_208[19:0];
  _RAND_209 = {1{`RANDOM}};
  tag_209 = _RAND_209[19:0];
  _RAND_210 = {1{`RANDOM}};
  tag_210 = _RAND_210[19:0];
  _RAND_211 = {1{`RANDOM}};
  tag_211 = _RAND_211[19:0];
  _RAND_212 = {1{`RANDOM}};
  tag_212 = _RAND_212[19:0];
  _RAND_213 = {1{`RANDOM}};
  tag_213 = _RAND_213[19:0];
  _RAND_214 = {1{`RANDOM}};
  tag_214 = _RAND_214[19:0];
  _RAND_215 = {1{`RANDOM}};
  tag_215 = _RAND_215[19:0];
  _RAND_216 = {1{`RANDOM}};
  tag_216 = _RAND_216[19:0];
  _RAND_217 = {1{`RANDOM}};
  tag_217 = _RAND_217[19:0];
  _RAND_218 = {1{`RANDOM}};
  tag_218 = _RAND_218[19:0];
  _RAND_219 = {1{`RANDOM}};
  tag_219 = _RAND_219[19:0];
  _RAND_220 = {1{`RANDOM}};
  tag_220 = _RAND_220[19:0];
  _RAND_221 = {1{`RANDOM}};
  tag_221 = _RAND_221[19:0];
  _RAND_222 = {1{`RANDOM}};
  tag_222 = _RAND_222[19:0];
  _RAND_223 = {1{`RANDOM}};
  tag_223 = _RAND_223[19:0];
  _RAND_224 = {1{`RANDOM}};
  tag_224 = _RAND_224[19:0];
  _RAND_225 = {1{`RANDOM}};
  tag_225 = _RAND_225[19:0];
  _RAND_226 = {1{`RANDOM}};
  tag_226 = _RAND_226[19:0];
  _RAND_227 = {1{`RANDOM}};
  tag_227 = _RAND_227[19:0];
  _RAND_228 = {1{`RANDOM}};
  tag_228 = _RAND_228[19:0];
  _RAND_229 = {1{`RANDOM}};
  tag_229 = _RAND_229[19:0];
  _RAND_230 = {1{`RANDOM}};
  tag_230 = _RAND_230[19:0];
  _RAND_231 = {1{`RANDOM}};
  tag_231 = _RAND_231[19:0];
  _RAND_232 = {1{`RANDOM}};
  tag_232 = _RAND_232[19:0];
  _RAND_233 = {1{`RANDOM}};
  tag_233 = _RAND_233[19:0];
  _RAND_234 = {1{`RANDOM}};
  tag_234 = _RAND_234[19:0];
  _RAND_235 = {1{`RANDOM}};
  tag_235 = _RAND_235[19:0];
  _RAND_236 = {1{`RANDOM}};
  tag_236 = _RAND_236[19:0];
  _RAND_237 = {1{`RANDOM}};
  tag_237 = _RAND_237[19:0];
  _RAND_238 = {1{`RANDOM}};
  tag_238 = _RAND_238[19:0];
  _RAND_239 = {1{`RANDOM}};
  tag_239 = _RAND_239[19:0];
  _RAND_240 = {1{`RANDOM}};
  tag_240 = _RAND_240[19:0];
  _RAND_241 = {1{`RANDOM}};
  tag_241 = _RAND_241[19:0];
  _RAND_242 = {1{`RANDOM}};
  tag_242 = _RAND_242[19:0];
  _RAND_243 = {1{`RANDOM}};
  tag_243 = _RAND_243[19:0];
  _RAND_244 = {1{`RANDOM}};
  tag_244 = _RAND_244[19:0];
  _RAND_245 = {1{`RANDOM}};
  tag_245 = _RAND_245[19:0];
  _RAND_246 = {1{`RANDOM}};
  tag_246 = _RAND_246[19:0];
  _RAND_247 = {1{`RANDOM}};
  tag_247 = _RAND_247[19:0];
  _RAND_248 = {1{`RANDOM}};
  tag_248 = _RAND_248[19:0];
  _RAND_249 = {1{`RANDOM}};
  tag_249 = _RAND_249[19:0];
  _RAND_250 = {1{`RANDOM}};
  tag_250 = _RAND_250[19:0];
  _RAND_251 = {1{`RANDOM}};
  tag_251 = _RAND_251[19:0];
  _RAND_252 = {1{`RANDOM}};
  tag_252 = _RAND_252[19:0];
  _RAND_253 = {1{`RANDOM}};
  tag_253 = _RAND_253[19:0];
  _RAND_254 = {1{`RANDOM}};
  tag_254 = _RAND_254[19:0];
  _RAND_255 = {1{`RANDOM}};
  tag_255 = _RAND_255[19:0];
  _RAND_256 = {1{`RANDOM}};
  valid_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_3 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_4 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_5 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_6 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_7 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_8 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_9 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_10 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_11 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_12 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_13 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_14 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_15 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_16 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_17 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_18 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_19 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_20 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_21 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_22 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_23 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_24 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_25 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_26 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_27 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_28 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_29 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_30 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_31 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_32 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_33 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_34 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_35 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_36 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_37 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_38 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_39 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_40 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_41 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_42 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_43 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_44 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_45 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_46 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_47 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_48 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_49 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_50 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_51 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_52 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_53 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_54 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_55 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_56 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_57 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_58 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_59 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_60 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_61 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_62 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_63 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_64 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_65 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_66 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_67 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid_68 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid_69 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid_70 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid_71 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid_72 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid_73 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid_74 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid_75 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid_76 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid_77 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid_78 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid_79 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid_80 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid_81 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid_82 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid_83 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid_84 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid_85 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid_86 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid_87 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid_88 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid_89 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid_90 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid_91 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid_92 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid_93 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid_94 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid_95 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid_96 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid_97 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid_98 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid_99 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid_100 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid_101 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid_102 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid_103 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid_104 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid_105 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid_106 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid_107 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid_108 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid_109 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid_110 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid_111 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid_112 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid_113 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid_114 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid_115 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid_116 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid_117 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid_118 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid_119 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid_120 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid_121 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid_122 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid_123 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid_124 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid_125 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid_126 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid_127 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  valid_128 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  valid_129 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  valid_130 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  valid_131 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  valid_132 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  valid_133 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  valid_134 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  valid_135 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  valid_136 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  valid_137 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  valid_138 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  valid_139 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  valid_140 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  valid_141 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  valid_142 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  valid_143 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  valid_144 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  valid_145 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  valid_146 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  valid_147 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  valid_148 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  valid_149 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  valid_150 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  valid_151 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  valid_152 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  valid_153 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  valid_154 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  valid_155 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  valid_156 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  valid_157 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  valid_158 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  valid_159 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  valid_160 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  valid_161 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  valid_162 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  valid_163 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  valid_164 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  valid_165 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  valid_166 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  valid_167 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  valid_168 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  valid_169 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  valid_170 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  valid_171 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  valid_172 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  valid_173 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  valid_174 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  valid_175 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  valid_176 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  valid_177 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  valid_178 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  valid_179 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  valid_180 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  valid_181 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  valid_182 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  valid_183 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  valid_184 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  valid_185 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  valid_186 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  valid_187 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  valid_188 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  valid_189 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  valid_190 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  valid_191 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  valid_192 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  valid_193 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  valid_194 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  valid_195 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  valid_196 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  valid_197 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  valid_198 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  valid_199 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  valid_200 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  valid_201 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  valid_202 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  valid_203 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  valid_204 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  valid_205 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  valid_206 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  valid_207 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  valid_208 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  valid_209 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  valid_210 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  valid_211 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  valid_212 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  valid_213 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  valid_214 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  valid_215 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  valid_216 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  valid_217 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  valid_218 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  valid_219 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  valid_220 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  valid_221 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  valid_222 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  valid_223 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  valid_224 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  valid_225 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  valid_226 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  valid_227 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  valid_228 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  valid_229 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  valid_230 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  valid_231 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  valid_232 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  valid_233 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  valid_234 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  valid_235 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  valid_236 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  valid_237 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  valid_238 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  valid_239 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  valid_240 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  valid_241 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  valid_242 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  valid_243 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  valid_244 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  valid_245 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  valid_246 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  valid_247 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  valid_248 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  valid_249 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  valid_250 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  valid_251 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  valid_252 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  valid_253 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  valid_254 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  valid_255 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  state = _RAND_512[1:0];
  _RAND_513 = {1{`RANDOM}};
  req_addr = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  cache_fill = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  cache_wen = _RAND_515[0:0];
  _RAND_516 = {4{`RANDOM}};
  cache_wdata = _RAND_516[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Dcache(
  input          clock,
  input          reset,
  input          io_dmem_data_valid,
  output         io_dmem_data_ready,
  input          io_dmem_data_req,
  input  [31:0]  io_dmem_data_addr,
  input  [1:0]   io_dmem_data_size,
  input  [7:0]   io_dmem_data_strb,
  output [63:0]  io_dmem_data_read,
  input  [63:0]  io_dmem_data_write,
  output         io_out_data_valid,
  input          io_out_data_ready,
  output         io_out_data_req,
  output [31:0]  io_out_data_addr,
  output [7:0]   io_out_data_strb,
  input  [127:0] io_out_data_read,
  output [127:0] io_out_data_write
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [127:0] _RAND_1028;
  reg [127:0] _RAND_1029;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] req_Q; // @[Dcache.scala 217:19]
  wire  req_CLK; // @[Dcache.scala 217:19]
  wire  req_CEN; // @[Dcache.scala 217:19]
  wire  req_WEN; // @[Dcache.scala 217:19]
  wire [127:0] req_BWEN; // @[Dcache.scala 217:19]
  wire [7:0] req_A; // @[Dcache.scala 217:19]
  wire [127:0] req_D; // @[Dcache.scala 217:19]
  reg [19:0] tag_0; // @[Dcache.scala 16:24]
  reg [19:0] tag_1; // @[Dcache.scala 16:24]
  reg [19:0] tag_2; // @[Dcache.scala 16:24]
  reg [19:0] tag_3; // @[Dcache.scala 16:24]
  reg [19:0] tag_4; // @[Dcache.scala 16:24]
  reg [19:0] tag_5; // @[Dcache.scala 16:24]
  reg [19:0] tag_6; // @[Dcache.scala 16:24]
  reg [19:0] tag_7; // @[Dcache.scala 16:24]
  reg [19:0] tag_8; // @[Dcache.scala 16:24]
  reg [19:0] tag_9; // @[Dcache.scala 16:24]
  reg [19:0] tag_10; // @[Dcache.scala 16:24]
  reg [19:0] tag_11; // @[Dcache.scala 16:24]
  reg [19:0] tag_12; // @[Dcache.scala 16:24]
  reg [19:0] tag_13; // @[Dcache.scala 16:24]
  reg [19:0] tag_14; // @[Dcache.scala 16:24]
  reg [19:0] tag_15; // @[Dcache.scala 16:24]
  reg [19:0] tag_16; // @[Dcache.scala 16:24]
  reg [19:0] tag_17; // @[Dcache.scala 16:24]
  reg [19:0] tag_18; // @[Dcache.scala 16:24]
  reg [19:0] tag_19; // @[Dcache.scala 16:24]
  reg [19:0] tag_20; // @[Dcache.scala 16:24]
  reg [19:0] tag_21; // @[Dcache.scala 16:24]
  reg [19:0] tag_22; // @[Dcache.scala 16:24]
  reg [19:0] tag_23; // @[Dcache.scala 16:24]
  reg [19:0] tag_24; // @[Dcache.scala 16:24]
  reg [19:0] tag_25; // @[Dcache.scala 16:24]
  reg [19:0] tag_26; // @[Dcache.scala 16:24]
  reg [19:0] tag_27; // @[Dcache.scala 16:24]
  reg [19:0] tag_28; // @[Dcache.scala 16:24]
  reg [19:0] tag_29; // @[Dcache.scala 16:24]
  reg [19:0] tag_30; // @[Dcache.scala 16:24]
  reg [19:0] tag_31; // @[Dcache.scala 16:24]
  reg [19:0] tag_32; // @[Dcache.scala 16:24]
  reg [19:0] tag_33; // @[Dcache.scala 16:24]
  reg [19:0] tag_34; // @[Dcache.scala 16:24]
  reg [19:0] tag_35; // @[Dcache.scala 16:24]
  reg [19:0] tag_36; // @[Dcache.scala 16:24]
  reg [19:0] tag_37; // @[Dcache.scala 16:24]
  reg [19:0] tag_38; // @[Dcache.scala 16:24]
  reg [19:0] tag_39; // @[Dcache.scala 16:24]
  reg [19:0] tag_40; // @[Dcache.scala 16:24]
  reg [19:0] tag_41; // @[Dcache.scala 16:24]
  reg [19:0] tag_42; // @[Dcache.scala 16:24]
  reg [19:0] tag_43; // @[Dcache.scala 16:24]
  reg [19:0] tag_44; // @[Dcache.scala 16:24]
  reg [19:0] tag_45; // @[Dcache.scala 16:24]
  reg [19:0] tag_46; // @[Dcache.scala 16:24]
  reg [19:0] tag_47; // @[Dcache.scala 16:24]
  reg [19:0] tag_48; // @[Dcache.scala 16:24]
  reg [19:0] tag_49; // @[Dcache.scala 16:24]
  reg [19:0] tag_50; // @[Dcache.scala 16:24]
  reg [19:0] tag_51; // @[Dcache.scala 16:24]
  reg [19:0] tag_52; // @[Dcache.scala 16:24]
  reg [19:0] tag_53; // @[Dcache.scala 16:24]
  reg [19:0] tag_54; // @[Dcache.scala 16:24]
  reg [19:0] tag_55; // @[Dcache.scala 16:24]
  reg [19:0] tag_56; // @[Dcache.scala 16:24]
  reg [19:0] tag_57; // @[Dcache.scala 16:24]
  reg [19:0] tag_58; // @[Dcache.scala 16:24]
  reg [19:0] tag_59; // @[Dcache.scala 16:24]
  reg [19:0] tag_60; // @[Dcache.scala 16:24]
  reg [19:0] tag_61; // @[Dcache.scala 16:24]
  reg [19:0] tag_62; // @[Dcache.scala 16:24]
  reg [19:0] tag_63; // @[Dcache.scala 16:24]
  reg [19:0] tag_64; // @[Dcache.scala 16:24]
  reg [19:0] tag_65; // @[Dcache.scala 16:24]
  reg [19:0] tag_66; // @[Dcache.scala 16:24]
  reg [19:0] tag_67; // @[Dcache.scala 16:24]
  reg [19:0] tag_68; // @[Dcache.scala 16:24]
  reg [19:0] tag_69; // @[Dcache.scala 16:24]
  reg [19:0] tag_70; // @[Dcache.scala 16:24]
  reg [19:0] tag_71; // @[Dcache.scala 16:24]
  reg [19:0] tag_72; // @[Dcache.scala 16:24]
  reg [19:0] tag_73; // @[Dcache.scala 16:24]
  reg [19:0] tag_74; // @[Dcache.scala 16:24]
  reg [19:0] tag_75; // @[Dcache.scala 16:24]
  reg [19:0] tag_76; // @[Dcache.scala 16:24]
  reg [19:0] tag_77; // @[Dcache.scala 16:24]
  reg [19:0] tag_78; // @[Dcache.scala 16:24]
  reg [19:0] tag_79; // @[Dcache.scala 16:24]
  reg [19:0] tag_80; // @[Dcache.scala 16:24]
  reg [19:0] tag_81; // @[Dcache.scala 16:24]
  reg [19:0] tag_82; // @[Dcache.scala 16:24]
  reg [19:0] tag_83; // @[Dcache.scala 16:24]
  reg [19:0] tag_84; // @[Dcache.scala 16:24]
  reg [19:0] tag_85; // @[Dcache.scala 16:24]
  reg [19:0] tag_86; // @[Dcache.scala 16:24]
  reg [19:0] tag_87; // @[Dcache.scala 16:24]
  reg [19:0] tag_88; // @[Dcache.scala 16:24]
  reg [19:0] tag_89; // @[Dcache.scala 16:24]
  reg [19:0] tag_90; // @[Dcache.scala 16:24]
  reg [19:0] tag_91; // @[Dcache.scala 16:24]
  reg [19:0] tag_92; // @[Dcache.scala 16:24]
  reg [19:0] tag_93; // @[Dcache.scala 16:24]
  reg [19:0] tag_94; // @[Dcache.scala 16:24]
  reg [19:0] tag_95; // @[Dcache.scala 16:24]
  reg [19:0] tag_96; // @[Dcache.scala 16:24]
  reg [19:0] tag_97; // @[Dcache.scala 16:24]
  reg [19:0] tag_98; // @[Dcache.scala 16:24]
  reg [19:0] tag_99; // @[Dcache.scala 16:24]
  reg [19:0] tag_100; // @[Dcache.scala 16:24]
  reg [19:0] tag_101; // @[Dcache.scala 16:24]
  reg [19:0] tag_102; // @[Dcache.scala 16:24]
  reg [19:0] tag_103; // @[Dcache.scala 16:24]
  reg [19:0] tag_104; // @[Dcache.scala 16:24]
  reg [19:0] tag_105; // @[Dcache.scala 16:24]
  reg [19:0] tag_106; // @[Dcache.scala 16:24]
  reg [19:0] tag_107; // @[Dcache.scala 16:24]
  reg [19:0] tag_108; // @[Dcache.scala 16:24]
  reg [19:0] tag_109; // @[Dcache.scala 16:24]
  reg [19:0] tag_110; // @[Dcache.scala 16:24]
  reg [19:0] tag_111; // @[Dcache.scala 16:24]
  reg [19:0] tag_112; // @[Dcache.scala 16:24]
  reg [19:0] tag_113; // @[Dcache.scala 16:24]
  reg [19:0] tag_114; // @[Dcache.scala 16:24]
  reg [19:0] tag_115; // @[Dcache.scala 16:24]
  reg [19:0] tag_116; // @[Dcache.scala 16:24]
  reg [19:0] tag_117; // @[Dcache.scala 16:24]
  reg [19:0] tag_118; // @[Dcache.scala 16:24]
  reg [19:0] tag_119; // @[Dcache.scala 16:24]
  reg [19:0] tag_120; // @[Dcache.scala 16:24]
  reg [19:0] tag_121; // @[Dcache.scala 16:24]
  reg [19:0] tag_122; // @[Dcache.scala 16:24]
  reg [19:0] tag_123; // @[Dcache.scala 16:24]
  reg [19:0] tag_124; // @[Dcache.scala 16:24]
  reg [19:0] tag_125; // @[Dcache.scala 16:24]
  reg [19:0] tag_126; // @[Dcache.scala 16:24]
  reg [19:0] tag_127; // @[Dcache.scala 16:24]
  reg [19:0] tag_128; // @[Dcache.scala 16:24]
  reg [19:0] tag_129; // @[Dcache.scala 16:24]
  reg [19:0] tag_130; // @[Dcache.scala 16:24]
  reg [19:0] tag_131; // @[Dcache.scala 16:24]
  reg [19:0] tag_132; // @[Dcache.scala 16:24]
  reg [19:0] tag_133; // @[Dcache.scala 16:24]
  reg [19:0] tag_134; // @[Dcache.scala 16:24]
  reg [19:0] tag_135; // @[Dcache.scala 16:24]
  reg [19:0] tag_136; // @[Dcache.scala 16:24]
  reg [19:0] tag_137; // @[Dcache.scala 16:24]
  reg [19:0] tag_138; // @[Dcache.scala 16:24]
  reg [19:0] tag_139; // @[Dcache.scala 16:24]
  reg [19:0] tag_140; // @[Dcache.scala 16:24]
  reg [19:0] tag_141; // @[Dcache.scala 16:24]
  reg [19:0] tag_142; // @[Dcache.scala 16:24]
  reg [19:0] tag_143; // @[Dcache.scala 16:24]
  reg [19:0] tag_144; // @[Dcache.scala 16:24]
  reg [19:0] tag_145; // @[Dcache.scala 16:24]
  reg [19:0] tag_146; // @[Dcache.scala 16:24]
  reg [19:0] tag_147; // @[Dcache.scala 16:24]
  reg [19:0] tag_148; // @[Dcache.scala 16:24]
  reg [19:0] tag_149; // @[Dcache.scala 16:24]
  reg [19:0] tag_150; // @[Dcache.scala 16:24]
  reg [19:0] tag_151; // @[Dcache.scala 16:24]
  reg [19:0] tag_152; // @[Dcache.scala 16:24]
  reg [19:0] tag_153; // @[Dcache.scala 16:24]
  reg [19:0] tag_154; // @[Dcache.scala 16:24]
  reg [19:0] tag_155; // @[Dcache.scala 16:24]
  reg [19:0] tag_156; // @[Dcache.scala 16:24]
  reg [19:0] tag_157; // @[Dcache.scala 16:24]
  reg [19:0] tag_158; // @[Dcache.scala 16:24]
  reg [19:0] tag_159; // @[Dcache.scala 16:24]
  reg [19:0] tag_160; // @[Dcache.scala 16:24]
  reg [19:0] tag_161; // @[Dcache.scala 16:24]
  reg [19:0] tag_162; // @[Dcache.scala 16:24]
  reg [19:0] tag_163; // @[Dcache.scala 16:24]
  reg [19:0] tag_164; // @[Dcache.scala 16:24]
  reg [19:0] tag_165; // @[Dcache.scala 16:24]
  reg [19:0] tag_166; // @[Dcache.scala 16:24]
  reg [19:0] tag_167; // @[Dcache.scala 16:24]
  reg [19:0] tag_168; // @[Dcache.scala 16:24]
  reg [19:0] tag_169; // @[Dcache.scala 16:24]
  reg [19:0] tag_170; // @[Dcache.scala 16:24]
  reg [19:0] tag_171; // @[Dcache.scala 16:24]
  reg [19:0] tag_172; // @[Dcache.scala 16:24]
  reg [19:0] tag_173; // @[Dcache.scala 16:24]
  reg [19:0] tag_174; // @[Dcache.scala 16:24]
  reg [19:0] tag_175; // @[Dcache.scala 16:24]
  reg [19:0] tag_176; // @[Dcache.scala 16:24]
  reg [19:0] tag_177; // @[Dcache.scala 16:24]
  reg [19:0] tag_178; // @[Dcache.scala 16:24]
  reg [19:0] tag_179; // @[Dcache.scala 16:24]
  reg [19:0] tag_180; // @[Dcache.scala 16:24]
  reg [19:0] tag_181; // @[Dcache.scala 16:24]
  reg [19:0] tag_182; // @[Dcache.scala 16:24]
  reg [19:0] tag_183; // @[Dcache.scala 16:24]
  reg [19:0] tag_184; // @[Dcache.scala 16:24]
  reg [19:0] tag_185; // @[Dcache.scala 16:24]
  reg [19:0] tag_186; // @[Dcache.scala 16:24]
  reg [19:0] tag_187; // @[Dcache.scala 16:24]
  reg [19:0] tag_188; // @[Dcache.scala 16:24]
  reg [19:0] tag_189; // @[Dcache.scala 16:24]
  reg [19:0] tag_190; // @[Dcache.scala 16:24]
  reg [19:0] tag_191; // @[Dcache.scala 16:24]
  reg [19:0] tag_192; // @[Dcache.scala 16:24]
  reg [19:0] tag_193; // @[Dcache.scala 16:24]
  reg [19:0] tag_194; // @[Dcache.scala 16:24]
  reg [19:0] tag_195; // @[Dcache.scala 16:24]
  reg [19:0] tag_196; // @[Dcache.scala 16:24]
  reg [19:0] tag_197; // @[Dcache.scala 16:24]
  reg [19:0] tag_198; // @[Dcache.scala 16:24]
  reg [19:0] tag_199; // @[Dcache.scala 16:24]
  reg [19:0] tag_200; // @[Dcache.scala 16:24]
  reg [19:0] tag_201; // @[Dcache.scala 16:24]
  reg [19:0] tag_202; // @[Dcache.scala 16:24]
  reg [19:0] tag_203; // @[Dcache.scala 16:24]
  reg [19:0] tag_204; // @[Dcache.scala 16:24]
  reg [19:0] tag_205; // @[Dcache.scala 16:24]
  reg [19:0] tag_206; // @[Dcache.scala 16:24]
  reg [19:0] tag_207; // @[Dcache.scala 16:24]
  reg [19:0] tag_208; // @[Dcache.scala 16:24]
  reg [19:0] tag_209; // @[Dcache.scala 16:24]
  reg [19:0] tag_210; // @[Dcache.scala 16:24]
  reg [19:0] tag_211; // @[Dcache.scala 16:24]
  reg [19:0] tag_212; // @[Dcache.scala 16:24]
  reg [19:0] tag_213; // @[Dcache.scala 16:24]
  reg [19:0] tag_214; // @[Dcache.scala 16:24]
  reg [19:0] tag_215; // @[Dcache.scala 16:24]
  reg [19:0] tag_216; // @[Dcache.scala 16:24]
  reg [19:0] tag_217; // @[Dcache.scala 16:24]
  reg [19:0] tag_218; // @[Dcache.scala 16:24]
  reg [19:0] tag_219; // @[Dcache.scala 16:24]
  reg [19:0] tag_220; // @[Dcache.scala 16:24]
  reg [19:0] tag_221; // @[Dcache.scala 16:24]
  reg [19:0] tag_222; // @[Dcache.scala 16:24]
  reg [19:0] tag_223; // @[Dcache.scala 16:24]
  reg [19:0] tag_224; // @[Dcache.scala 16:24]
  reg [19:0] tag_225; // @[Dcache.scala 16:24]
  reg [19:0] tag_226; // @[Dcache.scala 16:24]
  reg [19:0] tag_227; // @[Dcache.scala 16:24]
  reg [19:0] tag_228; // @[Dcache.scala 16:24]
  reg [19:0] tag_229; // @[Dcache.scala 16:24]
  reg [19:0] tag_230; // @[Dcache.scala 16:24]
  reg [19:0] tag_231; // @[Dcache.scala 16:24]
  reg [19:0] tag_232; // @[Dcache.scala 16:24]
  reg [19:0] tag_233; // @[Dcache.scala 16:24]
  reg [19:0] tag_234; // @[Dcache.scala 16:24]
  reg [19:0] tag_235; // @[Dcache.scala 16:24]
  reg [19:0] tag_236; // @[Dcache.scala 16:24]
  reg [19:0] tag_237; // @[Dcache.scala 16:24]
  reg [19:0] tag_238; // @[Dcache.scala 16:24]
  reg [19:0] tag_239; // @[Dcache.scala 16:24]
  reg [19:0] tag_240; // @[Dcache.scala 16:24]
  reg [19:0] tag_241; // @[Dcache.scala 16:24]
  reg [19:0] tag_242; // @[Dcache.scala 16:24]
  reg [19:0] tag_243; // @[Dcache.scala 16:24]
  reg [19:0] tag_244; // @[Dcache.scala 16:24]
  reg [19:0] tag_245; // @[Dcache.scala 16:24]
  reg [19:0] tag_246; // @[Dcache.scala 16:24]
  reg [19:0] tag_247; // @[Dcache.scala 16:24]
  reg [19:0] tag_248; // @[Dcache.scala 16:24]
  reg [19:0] tag_249; // @[Dcache.scala 16:24]
  reg [19:0] tag_250; // @[Dcache.scala 16:24]
  reg [19:0] tag_251; // @[Dcache.scala 16:24]
  reg [19:0] tag_252; // @[Dcache.scala 16:24]
  reg [19:0] tag_253; // @[Dcache.scala 16:24]
  reg [19:0] tag_254; // @[Dcache.scala 16:24]
  reg [19:0] tag_255; // @[Dcache.scala 16:24]
  reg  valid_0; // @[Dcache.scala 17:24]
  reg  valid_1; // @[Dcache.scala 17:24]
  reg  valid_2; // @[Dcache.scala 17:24]
  reg  valid_3; // @[Dcache.scala 17:24]
  reg  valid_4; // @[Dcache.scala 17:24]
  reg  valid_5; // @[Dcache.scala 17:24]
  reg  valid_6; // @[Dcache.scala 17:24]
  reg  valid_7; // @[Dcache.scala 17:24]
  reg  valid_8; // @[Dcache.scala 17:24]
  reg  valid_9; // @[Dcache.scala 17:24]
  reg  valid_10; // @[Dcache.scala 17:24]
  reg  valid_11; // @[Dcache.scala 17:24]
  reg  valid_12; // @[Dcache.scala 17:24]
  reg  valid_13; // @[Dcache.scala 17:24]
  reg  valid_14; // @[Dcache.scala 17:24]
  reg  valid_15; // @[Dcache.scala 17:24]
  reg  valid_16; // @[Dcache.scala 17:24]
  reg  valid_17; // @[Dcache.scala 17:24]
  reg  valid_18; // @[Dcache.scala 17:24]
  reg  valid_19; // @[Dcache.scala 17:24]
  reg  valid_20; // @[Dcache.scala 17:24]
  reg  valid_21; // @[Dcache.scala 17:24]
  reg  valid_22; // @[Dcache.scala 17:24]
  reg  valid_23; // @[Dcache.scala 17:24]
  reg  valid_24; // @[Dcache.scala 17:24]
  reg  valid_25; // @[Dcache.scala 17:24]
  reg  valid_26; // @[Dcache.scala 17:24]
  reg  valid_27; // @[Dcache.scala 17:24]
  reg  valid_28; // @[Dcache.scala 17:24]
  reg  valid_29; // @[Dcache.scala 17:24]
  reg  valid_30; // @[Dcache.scala 17:24]
  reg  valid_31; // @[Dcache.scala 17:24]
  reg  valid_32; // @[Dcache.scala 17:24]
  reg  valid_33; // @[Dcache.scala 17:24]
  reg  valid_34; // @[Dcache.scala 17:24]
  reg  valid_35; // @[Dcache.scala 17:24]
  reg  valid_36; // @[Dcache.scala 17:24]
  reg  valid_37; // @[Dcache.scala 17:24]
  reg  valid_38; // @[Dcache.scala 17:24]
  reg  valid_39; // @[Dcache.scala 17:24]
  reg  valid_40; // @[Dcache.scala 17:24]
  reg  valid_41; // @[Dcache.scala 17:24]
  reg  valid_42; // @[Dcache.scala 17:24]
  reg  valid_43; // @[Dcache.scala 17:24]
  reg  valid_44; // @[Dcache.scala 17:24]
  reg  valid_45; // @[Dcache.scala 17:24]
  reg  valid_46; // @[Dcache.scala 17:24]
  reg  valid_47; // @[Dcache.scala 17:24]
  reg  valid_48; // @[Dcache.scala 17:24]
  reg  valid_49; // @[Dcache.scala 17:24]
  reg  valid_50; // @[Dcache.scala 17:24]
  reg  valid_51; // @[Dcache.scala 17:24]
  reg  valid_52; // @[Dcache.scala 17:24]
  reg  valid_53; // @[Dcache.scala 17:24]
  reg  valid_54; // @[Dcache.scala 17:24]
  reg  valid_55; // @[Dcache.scala 17:24]
  reg  valid_56; // @[Dcache.scala 17:24]
  reg  valid_57; // @[Dcache.scala 17:24]
  reg  valid_58; // @[Dcache.scala 17:24]
  reg  valid_59; // @[Dcache.scala 17:24]
  reg  valid_60; // @[Dcache.scala 17:24]
  reg  valid_61; // @[Dcache.scala 17:24]
  reg  valid_62; // @[Dcache.scala 17:24]
  reg  valid_63; // @[Dcache.scala 17:24]
  reg  valid_64; // @[Dcache.scala 17:24]
  reg  valid_65; // @[Dcache.scala 17:24]
  reg  valid_66; // @[Dcache.scala 17:24]
  reg  valid_67; // @[Dcache.scala 17:24]
  reg  valid_68; // @[Dcache.scala 17:24]
  reg  valid_69; // @[Dcache.scala 17:24]
  reg  valid_70; // @[Dcache.scala 17:24]
  reg  valid_71; // @[Dcache.scala 17:24]
  reg  valid_72; // @[Dcache.scala 17:24]
  reg  valid_73; // @[Dcache.scala 17:24]
  reg  valid_74; // @[Dcache.scala 17:24]
  reg  valid_75; // @[Dcache.scala 17:24]
  reg  valid_76; // @[Dcache.scala 17:24]
  reg  valid_77; // @[Dcache.scala 17:24]
  reg  valid_78; // @[Dcache.scala 17:24]
  reg  valid_79; // @[Dcache.scala 17:24]
  reg  valid_80; // @[Dcache.scala 17:24]
  reg  valid_81; // @[Dcache.scala 17:24]
  reg  valid_82; // @[Dcache.scala 17:24]
  reg  valid_83; // @[Dcache.scala 17:24]
  reg  valid_84; // @[Dcache.scala 17:24]
  reg  valid_85; // @[Dcache.scala 17:24]
  reg  valid_86; // @[Dcache.scala 17:24]
  reg  valid_87; // @[Dcache.scala 17:24]
  reg  valid_88; // @[Dcache.scala 17:24]
  reg  valid_89; // @[Dcache.scala 17:24]
  reg  valid_90; // @[Dcache.scala 17:24]
  reg  valid_91; // @[Dcache.scala 17:24]
  reg  valid_92; // @[Dcache.scala 17:24]
  reg  valid_93; // @[Dcache.scala 17:24]
  reg  valid_94; // @[Dcache.scala 17:24]
  reg  valid_95; // @[Dcache.scala 17:24]
  reg  valid_96; // @[Dcache.scala 17:24]
  reg  valid_97; // @[Dcache.scala 17:24]
  reg  valid_98; // @[Dcache.scala 17:24]
  reg  valid_99; // @[Dcache.scala 17:24]
  reg  valid_100; // @[Dcache.scala 17:24]
  reg  valid_101; // @[Dcache.scala 17:24]
  reg  valid_102; // @[Dcache.scala 17:24]
  reg  valid_103; // @[Dcache.scala 17:24]
  reg  valid_104; // @[Dcache.scala 17:24]
  reg  valid_105; // @[Dcache.scala 17:24]
  reg  valid_106; // @[Dcache.scala 17:24]
  reg  valid_107; // @[Dcache.scala 17:24]
  reg  valid_108; // @[Dcache.scala 17:24]
  reg  valid_109; // @[Dcache.scala 17:24]
  reg  valid_110; // @[Dcache.scala 17:24]
  reg  valid_111; // @[Dcache.scala 17:24]
  reg  valid_112; // @[Dcache.scala 17:24]
  reg  valid_113; // @[Dcache.scala 17:24]
  reg  valid_114; // @[Dcache.scala 17:24]
  reg  valid_115; // @[Dcache.scala 17:24]
  reg  valid_116; // @[Dcache.scala 17:24]
  reg  valid_117; // @[Dcache.scala 17:24]
  reg  valid_118; // @[Dcache.scala 17:24]
  reg  valid_119; // @[Dcache.scala 17:24]
  reg  valid_120; // @[Dcache.scala 17:24]
  reg  valid_121; // @[Dcache.scala 17:24]
  reg  valid_122; // @[Dcache.scala 17:24]
  reg  valid_123; // @[Dcache.scala 17:24]
  reg  valid_124; // @[Dcache.scala 17:24]
  reg  valid_125; // @[Dcache.scala 17:24]
  reg  valid_126; // @[Dcache.scala 17:24]
  reg  valid_127; // @[Dcache.scala 17:24]
  reg  valid_128; // @[Dcache.scala 17:24]
  reg  valid_129; // @[Dcache.scala 17:24]
  reg  valid_130; // @[Dcache.scala 17:24]
  reg  valid_131; // @[Dcache.scala 17:24]
  reg  valid_132; // @[Dcache.scala 17:24]
  reg  valid_133; // @[Dcache.scala 17:24]
  reg  valid_134; // @[Dcache.scala 17:24]
  reg  valid_135; // @[Dcache.scala 17:24]
  reg  valid_136; // @[Dcache.scala 17:24]
  reg  valid_137; // @[Dcache.scala 17:24]
  reg  valid_138; // @[Dcache.scala 17:24]
  reg  valid_139; // @[Dcache.scala 17:24]
  reg  valid_140; // @[Dcache.scala 17:24]
  reg  valid_141; // @[Dcache.scala 17:24]
  reg  valid_142; // @[Dcache.scala 17:24]
  reg  valid_143; // @[Dcache.scala 17:24]
  reg  valid_144; // @[Dcache.scala 17:24]
  reg  valid_145; // @[Dcache.scala 17:24]
  reg  valid_146; // @[Dcache.scala 17:24]
  reg  valid_147; // @[Dcache.scala 17:24]
  reg  valid_148; // @[Dcache.scala 17:24]
  reg  valid_149; // @[Dcache.scala 17:24]
  reg  valid_150; // @[Dcache.scala 17:24]
  reg  valid_151; // @[Dcache.scala 17:24]
  reg  valid_152; // @[Dcache.scala 17:24]
  reg  valid_153; // @[Dcache.scala 17:24]
  reg  valid_154; // @[Dcache.scala 17:24]
  reg  valid_155; // @[Dcache.scala 17:24]
  reg  valid_156; // @[Dcache.scala 17:24]
  reg  valid_157; // @[Dcache.scala 17:24]
  reg  valid_158; // @[Dcache.scala 17:24]
  reg  valid_159; // @[Dcache.scala 17:24]
  reg  valid_160; // @[Dcache.scala 17:24]
  reg  valid_161; // @[Dcache.scala 17:24]
  reg  valid_162; // @[Dcache.scala 17:24]
  reg  valid_163; // @[Dcache.scala 17:24]
  reg  valid_164; // @[Dcache.scala 17:24]
  reg  valid_165; // @[Dcache.scala 17:24]
  reg  valid_166; // @[Dcache.scala 17:24]
  reg  valid_167; // @[Dcache.scala 17:24]
  reg  valid_168; // @[Dcache.scala 17:24]
  reg  valid_169; // @[Dcache.scala 17:24]
  reg  valid_170; // @[Dcache.scala 17:24]
  reg  valid_171; // @[Dcache.scala 17:24]
  reg  valid_172; // @[Dcache.scala 17:24]
  reg  valid_173; // @[Dcache.scala 17:24]
  reg  valid_174; // @[Dcache.scala 17:24]
  reg  valid_175; // @[Dcache.scala 17:24]
  reg  valid_176; // @[Dcache.scala 17:24]
  reg  valid_177; // @[Dcache.scala 17:24]
  reg  valid_178; // @[Dcache.scala 17:24]
  reg  valid_179; // @[Dcache.scala 17:24]
  reg  valid_180; // @[Dcache.scala 17:24]
  reg  valid_181; // @[Dcache.scala 17:24]
  reg  valid_182; // @[Dcache.scala 17:24]
  reg  valid_183; // @[Dcache.scala 17:24]
  reg  valid_184; // @[Dcache.scala 17:24]
  reg  valid_185; // @[Dcache.scala 17:24]
  reg  valid_186; // @[Dcache.scala 17:24]
  reg  valid_187; // @[Dcache.scala 17:24]
  reg  valid_188; // @[Dcache.scala 17:24]
  reg  valid_189; // @[Dcache.scala 17:24]
  reg  valid_190; // @[Dcache.scala 17:24]
  reg  valid_191; // @[Dcache.scala 17:24]
  reg  valid_192; // @[Dcache.scala 17:24]
  reg  valid_193; // @[Dcache.scala 17:24]
  reg  valid_194; // @[Dcache.scala 17:24]
  reg  valid_195; // @[Dcache.scala 17:24]
  reg  valid_196; // @[Dcache.scala 17:24]
  reg  valid_197; // @[Dcache.scala 17:24]
  reg  valid_198; // @[Dcache.scala 17:24]
  reg  valid_199; // @[Dcache.scala 17:24]
  reg  valid_200; // @[Dcache.scala 17:24]
  reg  valid_201; // @[Dcache.scala 17:24]
  reg  valid_202; // @[Dcache.scala 17:24]
  reg  valid_203; // @[Dcache.scala 17:24]
  reg  valid_204; // @[Dcache.scala 17:24]
  reg  valid_205; // @[Dcache.scala 17:24]
  reg  valid_206; // @[Dcache.scala 17:24]
  reg  valid_207; // @[Dcache.scala 17:24]
  reg  valid_208; // @[Dcache.scala 17:24]
  reg  valid_209; // @[Dcache.scala 17:24]
  reg  valid_210; // @[Dcache.scala 17:24]
  reg  valid_211; // @[Dcache.scala 17:24]
  reg  valid_212; // @[Dcache.scala 17:24]
  reg  valid_213; // @[Dcache.scala 17:24]
  reg  valid_214; // @[Dcache.scala 17:24]
  reg  valid_215; // @[Dcache.scala 17:24]
  reg  valid_216; // @[Dcache.scala 17:24]
  reg  valid_217; // @[Dcache.scala 17:24]
  reg  valid_218; // @[Dcache.scala 17:24]
  reg  valid_219; // @[Dcache.scala 17:24]
  reg  valid_220; // @[Dcache.scala 17:24]
  reg  valid_221; // @[Dcache.scala 17:24]
  reg  valid_222; // @[Dcache.scala 17:24]
  reg  valid_223; // @[Dcache.scala 17:24]
  reg  valid_224; // @[Dcache.scala 17:24]
  reg  valid_225; // @[Dcache.scala 17:24]
  reg  valid_226; // @[Dcache.scala 17:24]
  reg  valid_227; // @[Dcache.scala 17:24]
  reg  valid_228; // @[Dcache.scala 17:24]
  reg  valid_229; // @[Dcache.scala 17:24]
  reg  valid_230; // @[Dcache.scala 17:24]
  reg  valid_231; // @[Dcache.scala 17:24]
  reg  valid_232; // @[Dcache.scala 17:24]
  reg  valid_233; // @[Dcache.scala 17:24]
  reg  valid_234; // @[Dcache.scala 17:24]
  reg  valid_235; // @[Dcache.scala 17:24]
  reg  valid_236; // @[Dcache.scala 17:24]
  reg  valid_237; // @[Dcache.scala 17:24]
  reg  valid_238; // @[Dcache.scala 17:24]
  reg  valid_239; // @[Dcache.scala 17:24]
  reg  valid_240; // @[Dcache.scala 17:24]
  reg  valid_241; // @[Dcache.scala 17:24]
  reg  valid_242; // @[Dcache.scala 17:24]
  reg  valid_243; // @[Dcache.scala 17:24]
  reg  valid_244; // @[Dcache.scala 17:24]
  reg  valid_245; // @[Dcache.scala 17:24]
  reg  valid_246; // @[Dcache.scala 17:24]
  reg  valid_247; // @[Dcache.scala 17:24]
  reg  valid_248; // @[Dcache.scala 17:24]
  reg  valid_249; // @[Dcache.scala 17:24]
  reg  valid_250; // @[Dcache.scala 17:24]
  reg  valid_251; // @[Dcache.scala 17:24]
  reg  valid_252; // @[Dcache.scala 17:24]
  reg  valid_253; // @[Dcache.scala 17:24]
  reg  valid_254; // @[Dcache.scala 17:24]
  reg  valid_255; // @[Dcache.scala 17:24]
  reg  dirty_0; // @[Dcache.scala 18:24]
  reg  dirty_1; // @[Dcache.scala 18:24]
  reg  dirty_2; // @[Dcache.scala 18:24]
  reg  dirty_3; // @[Dcache.scala 18:24]
  reg  dirty_4; // @[Dcache.scala 18:24]
  reg  dirty_5; // @[Dcache.scala 18:24]
  reg  dirty_6; // @[Dcache.scala 18:24]
  reg  dirty_7; // @[Dcache.scala 18:24]
  reg  dirty_8; // @[Dcache.scala 18:24]
  reg  dirty_9; // @[Dcache.scala 18:24]
  reg  dirty_10; // @[Dcache.scala 18:24]
  reg  dirty_11; // @[Dcache.scala 18:24]
  reg  dirty_12; // @[Dcache.scala 18:24]
  reg  dirty_13; // @[Dcache.scala 18:24]
  reg  dirty_14; // @[Dcache.scala 18:24]
  reg  dirty_15; // @[Dcache.scala 18:24]
  reg  dirty_16; // @[Dcache.scala 18:24]
  reg  dirty_17; // @[Dcache.scala 18:24]
  reg  dirty_18; // @[Dcache.scala 18:24]
  reg  dirty_19; // @[Dcache.scala 18:24]
  reg  dirty_20; // @[Dcache.scala 18:24]
  reg  dirty_21; // @[Dcache.scala 18:24]
  reg  dirty_22; // @[Dcache.scala 18:24]
  reg  dirty_23; // @[Dcache.scala 18:24]
  reg  dirty_24; // @[Dcache.scala 18:24]
  reg  dirty_25; // @[Dcache.scala 18:24]
  reg  dirty_26; // @[Dcache.scala 18:24]
  reg  dirty_27; // @[Dcache.scala 18:24]
  reg  dirty_28; // @[Dcache.scala 18:24]
  reg  dirty_29; // @[Dcache.scala 18:24]
  reg  dirty_30; // @[Dcache.scala 18:24]
  reg  dirty_31; // @[Dcache.scala 18:24]
  reg  dirty_32; // @[Dcache.scala 18:24]
  reg  dirty_33; // @[Dcache.scala 18:24]
  reg  dirty_34; // @[Dcache.scala 18:24]
  reg  dirty_35; // @[Dcache.scala 18:24]
  reg  dirty_36; // @[Dcache.scala 18:24]
  reg  dirty_37; // @[Dcache.scala 18:24]
  reg  dirty_38; // @[Dcache.scala 18:24]
  reg  dirty_39; // @[Dcache.scala 18:24]
  reg  dirty_40; // @[Dcache.scala 18:24]
  reg  dirty_41; // @[Dcache.scala 18:24]
  reg  dirty_42; // @[Dcache.scala 18:24]
  reg  dirty_43; // @[Dcache.scala 18:24]
  reg  dirty_44; // @[Dcache.scala 18:24]
  reg  dirty_45; // @[Dcache.scala 18:24]
  reg  dirty_46; // @[Dcache.scala 18:24]
  reg  dirty_47; // @[Dcache.scala 18:24]
  reg  dirty_48; // @[Dcache.scala 18:24]
  reg  dirty_49; // @[Dcache.scala 18:24]
  reg  dirty_50; // @[Dcache.scala 18:24]
  reg  dirty_51; // @[Dcache.scala 18:24]
  reg  dirty_52; // @[Dcache.scala 18:24]
  reg  dirty_53; // @[Dcache.scala 18:24]
  reg  dirty_54; // @[Dcache.scala 18:24]
  reg  dirty_55; // @[Dcache.scala 18:24]
  reg  dirty_56; // @[Dcache.scala 18:24]
  reg  dirty_57; // @[Dcache.scala 18:24]
  reg  dirty_58; // @[Dcache.scala 18:24]
  reg  dirty_59; // @[Dcache.scala 18:24]
  reg  dirty_60; // @[Dcache.scala 18:24]
  reg  dirty_61; // @[Dcache.scala 18:24]
  reg  dirty_62; // @[Dcache.scala 18:24]
  reg  dirty_63; // @[Dcache.scala 18:24]
  reg  dirty_64; // @[Dcache.scala 18:24]
  reg  dirty_65; // @[Dcache.scala 18:24]
  reg  dirty_66; // @[Dcache.scala 18:24]
  reg  dirty_67; // @[Dcache.scala 18:24]
  reg  dirty_68; // @[Dcache.scala 18:24]
  reg  dirty_69; // @[Dcache.scala 18:24]
  reg  dirty_70; // @[Dcache.scala 18:24]
  reg  dirty_71; // @[Dcache.scala 18:24]
  reg  dirty_72; // @[Dcache.scala 18:24]
  reg  dirty_73; // @[Dcache.scala 18:24]
  reg  dirty_74; // @[Dcache.scala 18:24]
  reg  dirty_75; // @[Dcache.scala 18:24]
  reg  dirty_76; // @[Dcache.scala 18:24]
  reg  dirty_77; // @[Dcache.scala 18:24]
  reg  dirty_78; // @[Dcache.scala 18:24]
  reg  dirty_79; // @[Dcache.scala 18:24]
  reg  dirty_80; // @[Dcache.scala 18:24]
  reg  dirty_81; // @[Dcache.scala 18:24]
  reg  dirty_82; // @[Dcache.scala 18:24]
  reg  dirty_83; // @[Dcache.scala 18:24]
  reg  dirty_84; // @[Dcache.scala 18:24]
  reg  dirty_85; // @[Dcache.scala 18:24]
  reg  dirty_86; // @[Dcache.scala 18:24]
  reg  dirty_87; // @[Dcache.scala 18:24]
  reg  dirty_88; // @[Dcache.scala 18:24]
  reg  dirty_89; // @[Dcache.scala 18:24]
  reg  dirty_90; // @[Dcache.scala 18:24]
  reg  dirty_91; // @[Dcache.scala 18:24]
  reg  dirty_92; // @[Dcache.scala 18:24]
  reg  dirty_93; // @[Dcache.scala 18:24]
  reg  dirty_94; // @[Dcache.scala 18:24]
  reg  dirty_95; // @[Dcache.scala 18:24]
  reg  dirty_96; // @[Dcache.scala 18:24]
  reg  dirty_97; // @[Dcache.scala 18:24]
  reg  dirty_98; // @[Dcache.scala 18:24]
  reg  dirty_99; // @[Dcache.scala 18:24]
  reg  dirty_100; // @[Dcache.scala 18:24]
  reg  dirty_101; // @[Dcache.scala 18:24]
  reg  dirty_102; // @[Dcache.scala 18:24]
  reg  dirty_103; // @[Dcache.scala 18:24]
  reg  dirty_104; // @[Dcache.scala 18:24]
  reg  dirty_105; // @[Dcache.scala 18:24]
  reg  dirty_106; // @[Dcache.scala 18:24]
  reg  dirty_107; // @[Dcache.scala 18:24]
  reg  dirty_108; // @[Dcache.scala 18:24]
  reg  dirty_109; // @[Dcache.scala 18:24]
  reg  dirty_110; // @[Dcache.scala 18:24]
  reg  dirty_111; // @[Dcache.scala 18:24]
  reg  dirty_112; // @[Dcache.scala 18:24]
  reg  dirty_113; // @[Dcache.scala 18:24]
  reg  dirty_114; // @[Dcache.scala 18:24]
  reg  dirty_115; // @[Dcache.scala 18:24]
  reg  dirty_116; // @[Dcache.scala 18:24]
  reg  dirty_117; // @[Dcache.scala 18:24]
  reg  dirty_118; // @[Dcache.scala 18:24]
  reg  dirty_119; // @[Dcache.scala 18:24]
  reg  dirty_120; // @[Dcache.scala 18:24]
  reg  dirty_121; // @[Dcache.scala 18:24]
  reg  dirty_122; // @[Dcache.scala 18:24]
  reg  dirty_123; // @[Dcache.scala 18:24]
  reg  dirty_124; // @[Dcache.scala 18:24]
  reg  dirty_125; // @[Dcache.scala 18:24]
  reg  dirty_126; // @[Dcache.scala 18:24]
  reg  dirty_127; // @[Dcache.scala 18:24]
  reg  dirty_128; // @[Dcache.scala 18:24]
  reg  dirty_129; // @[Dcache.scala 18:24]
  reg  dirty_130; // @[Dcache.scala 18:24]
  reg  dirty_131; // @[Dcache.scala 18:24]
  reg  dirty_132; // @[Dcache.scala 18:24]
  reg  dirty_133; // @[Dcache.scala 18:24]
  reg  dirty_134; // @[Dcache.scala 18:24]
  reg  dirty_135; // @[Dcache.scala 18:24]
  reg  dirty_136; // @[Dcache.scala 18:24]
  reg  dirty_137; // @[Dcache.scala 18:24]
  reg  dirty_138; // @[Dcache.scala 18:24]
  reg  dirty_139; // @[Dcache.scala 18:24]
  reg  dirty_140; // @[Dcache.scala 18:24]
  reg  dirty_141; // @[Dcache.scala 18:24]
  reg  dirty_142; // @[Dcache.scala 18:24]
  reg  dirty_143; // @[Dcache.scala 18:24]
  reg  dirty_144; // @[Dcache.scala 18:24]
  reg  dirty_145; // @[Dcache.scala 18:24]
  reg  dirty_146; // @[Dcache.scala 18:24]
  reg  dirty_147; // @[Dcache.scala 18:24]
  reg  dirty_148; // @[Dcache.scala 18:24]
  reg  dirty_149; // @[Dcache.scala 18:24]
  reg  dirty_150; // @[Dcache.scala 18:24]
  reg  dirty_151; // @[Dcache.scala 18:24]
  reg  dirty_152; // @[Dcache.scala 18:24]
  reg  dirty_153; // @[Dcache.scala 18:24]
  reg  dirty_154; // @[Dcache.scala 18:24]
  reg  dirty_155; // @[Dcache.scala 18:24]
  reg  dirty_156; // @[Dcache.scala 18:24]
  reg  dirty_157; // @[Dcache.scala 18:24]
  reg  dirty_158; // @[Dcache.scala 18:24]
  reg  dirty_159; // @[Dcache.scala 18:24]
  reg  dirty_160; // @[Dcache.scala 18:24]
  reg  dirty_161; // @[Dcache.scala 18:24]
  reg  dirty_162; // @[Dcache.scala 18:24]
  reg  dirty_163; // @[Dcache.scala 18:24]
  reg  dirty_164; // @[Dcache.scala 18:24]
  reg  dirty_165; // @[Dcache.scala 18:24]
  reg  dirty_166; // @[Dcache.scala 18:24]
  reg  dirty_167; // @[Dcache.scala 18:24]
  reg  dirty_168; // @[Dcache.scala 18:24]
  reg  dirty_169; // @[Dcache.scala 18:24]
  reg  dirty_170; // @[Dcache.scala 18:24]
  reg  dirty_171; // @[Dcache.scala 18:24]
  reg  dirty_172; // @[Dcache.scala 18:24]
  reg  dirty_173; // @[Dcache.scala 18:24]
  reg  dirty_174; // @[Dcache.scala 18:24]
  reg  dirty_175; // @[Dcache.scala 18:24]
  reg  dirty_176; // @[Dcache.scala 18:24]
  reg  dirty_177; // @[Dcache.scala 18:24]
  reg  dirty_178; // @[Dcache.scala 18:24]
  reg  dirty_179; // @[Dcache.scala 18:24]
  reg  dirty_180; // @[Dcache.scala 18:24]
  reg  dirty_181; // @[Dcache.scala 18:24]
  reg  dirty_182; // @[Dcache.scala 18:24]
  reg  dirty_183; // @[Dcache.scala 18:24]
  reg  dirty_184; // @[Dcache.scala 18:24]
  reg  dirty_185; // @[Dcache.scala 18:24]
  reg  dirty_186; // @[Dcache.scala 18:24]
  reg  dirty_187; // @[Dcache.scala 18:24]
  reg  dirty_188; // @[Dcache.scala 18:24]
  reg  dirty_189; // @[Dcache.scala 18:24]
  reg  dirty_190; // @[Dcache.scala 18:24]
  reg  dirty_191; // @[Dcache.scala 18:24]
  reg  dirty_192; // @[Dcache.scala 18:24]
  reg  dirty_193; // @[Dcache.scala 18:24]
  reg  dirty_194; // @[Dcache.scala 18:24]
  reg  dirty_195; // @[Dcache.scala 18:24]
  reg  dirty_196; // @[Dcache.scala 18:24]
  reg  dirty_197; // @[Dcache.scala 18:24]
  reg  dirty_198; // @[Dcache.scala 18:24]
  reg  dirty_199; // @[Dcache.scala 18:24]
  reg  dirty_200; // @[Dcache.scala 18:24]
  reg  dirty_201; // @[Dcache.scala 18:24]
  reg  dirty_202; // @[Dcache.scala 18:24]
  reg  dirty_203; // @[Dcache.scala 18:24]
  reg  dirty_204; // @[Dcache.scala 18:24]
  reg  dirty_205; // @[Dcache.scala 18:24]
  reg  dirty_206; // @[Dcache.scala 18:24]
  reg  dirty_207; // @[Dcache.scala 18:24]
  reg  dirty_208; // @[Dcache.scala 18:24]
  reg  dirty_209; // @[Dcache.scala 18:24]
  reg  dirty_210; // @[Dcache.scala 18:24]
  reg  dirty_211; // @[Dcache.scala 18:24]
  reg  dirty_212; // @[Dcache.scala 18:24]
  reg  dirty_213; // @[Dcache.scala 18:24]
  reg  dirty_214; // @[Dcache.scala 18:24]
  reg  dirty_215; // @[Dcache.scala 18:24]
  reg  dirty_216; // @[Dcache.scala 18:24]
  reg  dirty_217; // @[Dcache.scala 18:24]
  reg  dirty_218; // @[Dcache.scala 18:24]
  reg  dirty_219; // @[Dcache.scala 18:24]
  reg  dirty_220; // @[Dcache.scala 18:24]
  reg  dirty_221; // @[Dcache.scala 18:24]
  reg  dirty_222; // @[Dcache.scala 18:24]
  reg  dirty_223; // @[Dcache.scala 18:24]
  reg  dirty_224; // @[Dcache.scala 18:24]
  reg  dirty_225; // @[Dcache.scala 18:24]
  reg  dirty_226; // @[Dcache.scala 18:24]
  reg  dirty_227; // @[Dcache.scala 18:24]
  reg  dirty_228; // @[Dcache.scala 18:24]
  reg  dirty_229; // @[Dcache.scala 18:24]
  reg  dirty_230; // @[Dcache.scala 18:24]
  reg  dirty_231; // @[Dcache.scala 18:24]
  reg  dirty_232; // @[Dcache.scala 18:24]
  reg  dirty_233; // @[Dcache.scala 18:24]
  reg  dirty_234; // @[Dcache.scala 18:24]
  reg  dirty_235; // @[Dcache.scala 18:24]
  reg  dirty_236; // @[Dcache.scala 18:24]
  reg  dirty_237; // @[Dcache.scala 18:24]
  reg  dirty_238; // @[Dcache.scala 18:24]
  reg  dirty_239; // @[Dcache.scala 18:24]
  reg  dirty_240; // @[Dcache.scala 18:24]
  reg  dirty_241; // @[Dcache.scala 18:24]
  reg  dirty_242; // @[Dcache.scala 18:24]
  reg  dirty_243; // @[Dcache.scala 18:24]
  reg  dirty_244; // @[Dcache.scala 18:24]
  reg  dirty_245; // @[Dcache.scala 18:24]
  reg  dirty_246; // @[Dcache.scala 18:24]
  reg  dirty_247; // @[Dcache.scala 18:24]
  reg  dirty_248; // @[Dcache.scala 18:24]
  reg  dirty_249; // @[Dcache.scala 18:24]
  reg  dirty_250; // @[Dcache.scala 18:24]
  reg  dirty_251; // @[Dcache.scala 18:24]
  reg  dirty_252; // @[Dcache.scala 18:24]
  reg  dirty_253; // @[Dcache.scala 18:24]
  reg  dirty_254; // @[Dcache.scala 18:24]
  reg  dirty_255; // @[Dcache.scala 18:24]
  reg [3:0] offset_0; // @[Dcache.scala 19:24]
  reg [3:0] offset_1; // @[Dcache.scala 19:24]
  reg [3:0] offset_2; // @[Dcache.scala 19:24]
  reg [3:0] offset_3; // @[Dcache.scala 19:24]
  reg [3:0] offset_4; // @[Dcache.scala 19:24]
  reg [3:0] offset_5; // @[Dcache.scala 19:24]
  reg [3:0] offset_6; // @[Dcache.scala 19:24]
  reg [3:0] offset_7; // @[Dcache.scala 19:24]
  reg [3:0] offset_8; // @[Dcache.scala 19:24]
  reg [3:0] offset_9; // @[Dcache.scala 19:24]
  reg [3:0] offset_10; // @[Dcache.scala 19:24]
  reg [3:0] offset_11; // @[Dcache.scala 19:24]
  reg [3:0] offset_12; // @[Dcache.scala 19:24]
  reg [3:0] offset_13; // @[Dcache.scala 19:24]
  reg [3:0] offset_14; // @[Dcache.scala 19:24]
  reg [3:0] offset_15; // @[Dcache.scala 19:24]
  reg [3:0] offset_16; // @[Dcache.scala 19:24]
  reg [3:0] offset_17; // @[Dcache.scala 19:24]
  reg [3:0] offset_18; // @[Dcache.scala 19:24]
  reg [3:0] offset_19; // @[Dcache.scala 19:24]
  reg [3:0] offset_20; // @[Dcache.scala 19:24]
  reg [3:0] offset_21; // @[Dcache.scala 19:24]
  reg [3:0] offset_22; // @[Dcache.scala 19:24]
  reg [3:0] offset_23; // @[Dcache.scala 19:24]
  reg [3:0] offset_24; // @[Dcache.scala 19:24]
  reg [3:0] offset_25; // @[Dcache.scala 19:24]
  reg [3:0] offset_26; // @[Dcache.scala 19:24]
  reg [3:0] offset_27; // @[Dcache.scala 19:24]
  reg [3:0] offset_28; // @[Dcache.scala 19:24]
  reg [3:0] offset_29; // @[Dcache.scala 19:24]
  reg [3:0] offset_30; // @[Dcache.scala 19:24]
  reg [3:0] offset_31; // @[Dcache.scala 19:24]
  reg [3:0] offset_32; // @[Dcache.scala 19:24]
  reg [3:0] offset_33; // @[Dcache.scala 19:24]
  reg [3:0] offset_34; // @[Dcache.scala 19:24]
  reg [3:0] offset_35; // @[Dcache.scala 19:24]
  reg [3:0] offset_36; // @[Dcache.scala 19:24]
  reg [3:0] offset_37; // @[Dcache.scala 19:24]
  reg [3:0] offset_38; // @[Dcache.scala 19:24]
  reg [3:0] offset_39; // @[Dcache.scala 19:24]
  reg [3:0] offset_40; // @[Dcache.scala 19:24]
  reg [3:0] offset_41; // @[Dcache.scala 19:24]
  reg [3:0] offset_42; // @[Dcache.scala 19:24]
  reg [3:0] offset_43; // @[Dcache.scala 19:24]
  reg [3:0] offset_44; // @[Dcache.scala 19:24]
  reg [3:0] offset_45; // @[Dcache.scala 19:24]
  reg [3:0] offset_46; // @[Dcache.scala 19:24]
  reg [3:0] offset_47; // @[Dcache.scala 19:24]
  reg [3:0] offset_48; // @[Dcache.scala 19:24]
  reg [3:0] offset_49; // @[Dcache.scala 19:24]
  reg [3:0] offset_50; // @[Dcache.scala 19:24]
  reg [3:0] offset_51; // @[Dcache.scala 19:24]
  reg [3:0] offset_52; // @[Dcache.scala 19:24]
  reg [3:0] offset_53; // @[Dcache.scala 19:24]
  reg [3:0] offset_54; // @[Dcache.scala 19:24]
  reg [3:0] offset_55; // @[Dcache.scala 19:24]
  reg [3:0] offset_56; // @[Dcache.scala 19:24]
  reg [3:0] offset_57; // @[Dcache.scala 19:24]
  reg [3:0] offset_58; // @[Dcache.scala 19:24]
  reg [3:0] offset_59; // @[Dcache.scala 19:24]
  reg [3:0] offset_60; // @[Dcache.scala 19:24]
  reg [3:0] offset_61; // @[Dcache.scala 19:24]
  reg [3:0] offset_62; // @[Dcache.scala 19:24]
  reg [3:0] offset_63; // @[Dcache.scala 19:24]
  reg [3:0] offset_64; // @[Dcache.scala 19:24]
  reg [3:0] offset_65; // @[Dcache.scala 19:24]
  reg [3:0] offset_66; // @[Dcache.scala 19:24]
  reg [3:0] offset_67; // @[Dcache.scala 19:24]
  reg [3:0] offset_68; // @[Dcache.scala 19:24]
  reg [3:0] offset_69; // @[Dcache.scala 19:24]
  reg [3:0] offset_70; // @[Dcache.scala 19:24]
  reg [3:0] offset_71; // @[Dcache.scala 19:24]
  reg [3:0] offset_72; // @[Dcache.scala 19:24]
  reg [3:0] offset_73; // @[Dcache.scala 19:24]
  reg [3:0] offset_74; // @[Dcache.scala 19:24]
  reg [3:0] offset_75; // @[Dcache.scala 19:24]
  reg [3:0] offset_76; // @[Dcache.scala 19:24]
  reg [3:0] offset_77; // @[Dcache.scala 19:24]
  reg [3:0] offset_78; // @[Dcache.scala 19:24]
  reg [3:0] offset_79; // @[Dcache.scala 19:24]
  reg [3:0] offset_80; // @[Dcache.scala 19:24]
  reg [3:0] offset_81; // @[Dcache.scala 19:24]
  reg [3:0] offset_82; // @[Dcache.scala 19:24]
  reg [3:0] offset_83; // @[Dcache.scala 19:24]
  reg [3:0] offset_84; // @[Dcache.scala 19:24]
  reg [3:0] offset_85; // @[Dcache.scala 19:24]
  reg [3:0] offset_86; // @[Dcache.scala 19:24]
  reg [3:0] offset_87; // @[Dcache.scala 19:24]
  reg [3:0] offset_88; // @[Dcache.scala 19:24]
  reg [3:0] offset_89; // @[Dcache.scala 19:24]
  reg [3:0] offset_90; // @[Dcache.scala 19:24]
  reg [3:0] offset_91; // @[Dcache.scala 19:24]
  reg [3:0] offset_92; // @[Dcache.scala 19:24]
  reg [3:0] offset_93; // @[Dcache.scala 19:24]
  reg [3:0] offset_94; // @[Dcache.scala 19:24]
  reg [3:0] offset_95; // @[Dcache.scala 19:24]
  reg [3:0] offset_96; // @[Dcache.scala 19:24]
  reg [3:0] offset_97; // @[Dcache.scala 19:24]
  reg [3:0] offset_98; // @[Dcache.scala 19:24]
  reg [3:0] offset_99; // @[Dcache.scala 19:24]
  reg [3:0] offset_100; // @[Dcache.scala 19:24]
  reg [3:0] offset_101; // @[Dcache.scala 19:24]
  reg [3:0] offset_102; // @[Dcache.scala 19:24]
  reg [3:0] offset_103; // @[Dcache.scala 19:24]
  reg [3:0] offset_104; // @[Dcache.scala 19:24]
  reg [3:0] offset_105; // @[Dcache.scala 19:24]
  reg [3:0] offset_106; // @[Dcache.scala 19:24]
  reg [3:0] offset_107; // @[Dcache.scala 19:24]
  reg [3:0] offset_108; // @[Dcache.scala 19:24]
  reg [3:0] offset_109; // @[Dcache.scala 19:24]
  reg [3:0] offset_110; // @[Dcache.scala 19:24]
  reg [3:0] offset_111; // @[Dcache.scala 19:24]
  reg [3:0] offset_112; // @[Dcache.scala 19:24]
  reg [3:0] offset_113; // @[Dcache.scala 19:24]
  reg [3:0] offset_114; // @[Dcache.scala 19:24]
  reg [3:0] offset_115; // @[Dcache.scala 19:24]
  reg [3:0] offset_116; // @[Dcache.scala 19:24]
  reg [3:0] offset_117; // @[Dcache.scala 19:24]
  reg [3:0] offset_118; // @[Dcache.scala 19:24]
  reg [3:0] offset_119; // @[Dcache.scala 19:24]
  reg [3:0] offset_120; // @[Dcache.scala 19:24]
  reg [3:0] offset_121; // @[Dcache.scala 19:24]
  reg [3:0] offset_122; // @[Dcache.scala 19:24]
  reg [3:0] offset_123; // @[Dcache.scala 19:24]
  reg [3:0] offset_124; // @[Dcache.scala 19:24]
  reg [3:0] offset_125; // @[Dcache.scala 19:24]
  reg [3:0] offset_126; // @[Dcache.scala 19:24]
  reg [3:0] offset_127; // @[Dcache.scala 19:24]
  reg [3:0] offset_128; // @[Dcache.scala 19:24]
  reg [3:0] offset_129; // @[Dcache.scala 19:24]
  reg [3:0] offset_130; // @[Dcache.scala 19:24]
  reg [3:0] offset_131; // @[Dcache.scala 19:24]
  reg [3:0] offset_132; // @[Dcache.scala 19:24]
  reg [3:0] offset_133; // @[Dcache.scala 19:24]
  reg [3:0] offset_134; // @[Dcache.scala 19:24]
  reg [3:0] offset_135; // @[Dcache.scala 19:24]
  reg [3:0] offset_136; // @[Dcache.scala 19:24]
  reg [3:0] offset_137; // @[Dcache.scala 19:24]
  reg [3:0] offset_138; // @[Dcache.scala 19:24]
  reg [3:0] offset_139; // @[Dcache.scala 19:24]
  reg [3:0] offset_140; // @[Dcache.scala 19:24]
  reg [3:0] offset_141; // @[Dcache.scala 19:24]
  reg [3:0] offset_142; // @[Dcache.scala 19:24]
  reg [3:0] offset_143; // @[Dcache.scala 19:24]
  reg [3:0] offset_144; // @[Dcache.scala 19:24]
  reg [3:0] offset_145; // @[Dcache.scala 19:24]
  reg [3:0] offset_146; // @[Dcache.scala 19:24]
  reg [3:0] offset_147; // @[Dcache.scala 19:24]
  reg [3:0] offset_148; // @[Dcache.scala 19:24]
  reg [3:0] offset_149; // @[Dcache.scala 19:24]
  reg [3:0] offset_150; // @[Dcache.scala 19:24]
  reg [3:0] offset_151; // @[Dcache.scala 19:24]
  reg [3:0] offset_152; // @[Dcache.scala 19:24]
  reg [3:0] offset_153; // @[Dcache.scala 19:24]
  reg [3:0] offset_154; // @[Dcache.scala 19:24]
  reg [3:0] offset_155; // @[Dcache.scala 19:24]
  reg [3:0] offset_156; // @[Dcache.scala 19:24]
  reg [3:0] offset_157; // @[Dcache.scala 19:24]
  reg [3:0] offset_158; // @[Dcache.scala 19:24]
  reg [3:0] offset_159; // @[Dcache.scala 19:24]
  reg [3:0] offset_160; // @[Dcache.scala 19:24]
  reg [3:0] offset_161; // @[Dcache.scala 19:24]
  reg [3:0] offset_162; // @[Dcache.scala 19:24]
  reg [3:0] offset_163; // @[Dcache.scala 19:24]
  reg [3:0] offset_164; // @[Dcache.scala 19:24]
  reg [3:0] offset_165; // @[Dcache.scala 19:24]
  reg [3:0] offset_166; // @[Dcache.scala 19:24]
  reg [3:0] offset_167; // @[Dcache.scala 19:24]
  reg [3:0] offset_168; // @[Dcache.scala 19:24]
  reg [3:0] offset_169; // @[Dcache.scala 19:24]
  reg [3:0] offset_170; // @[Dcache.scala 19:24]
  reg [3:0] offset_171; // @[Dcache.scala 19:24]
  reg [3:0] offset_172; // @[Dcache.scala 19:24]
  reg [3:0] offset_173; // @[Dcache.scala 19:24]
  reg [3:0] offset_174; // @[Dcache.scala 19:24]
  reg [3:0] offset_175; // @[Dcache.scala 19:24]
  reg [3:0] offset_176; // @[Dcache.scala 19:24]
  reg [3:0] offset_177; // @[Dcache.scala 19:24]
  reg [3:0] offset_178; // @[Dcache.scala 19:24]
  reg [3:0] offset_179; // @[Dcache.scala 19:24]
  reg [3:0] offset_180; // @[Dcache.scala 19:24]
  reg [3:0] offset_181; // @[Dcache.scala 19:24]
  reg [3:0] offset_182; // @[Dcache.scala 19:24]
  reg [3:0] offset_183; // @[Dcache.scala 19:24]
  reg [3:0] offset_184; // @[Dcache.scala 19:24]
  reg [3:0] offset_185; // @[Dcache.scala 19:24]
  reg [3:0] offset_186; // @[Dcache.scala 19:24]
  reg [3:0] offset_187; // @[Dcache.scala 19:24]
  reg [3:0] offset_188; // @[Dcache.scala 19:24]
  reg [3:0] offset_189; // @[Dcache.scala 19:24]
  reg [3:0] offset_190; // @[Dcache.scala 19:24]
  reg [3:0] offset_191; // @[Dcache.scala 19:24]
  reg [3:0] offset_192; // @[Dcache.scala 19:24]
  reg [3:0] offset_193; // @[Dcache.scala 19:24]
  reg [3:0] offset_194; // @[Dcache.scala 19:24]
  reg [3:0] offset_195; // @[Dcache.scala 19:24]
  reg [3:0] offset_196; // @[Dcache.scala 19:24]
  reg [3:0] offset_197; // @[Dcache.scala 19:24]
  reg [3:0] offset_198; // @[Dcache.scala 19:24]
  reg [3:0] offset_199; // @[Dcache.scala 19:24]
  reg [3:0] offset_200; // @[Dcache.scala 19:24]
  reg [3:0] offset_201; // @[Dcache.scala 19:24]
  reg [3:0] offset_202; // @[Dcache.scala 19:24]
  reg [3:0] offset_203; // @[Dcache.scala 19:24]
  reg [3:0] offset_204; // @[Dcache.scala 19:24]
  reg [3:0] offset_205; // @[Dcache.scala 19:24]
  reg [3:0] offset_206; // @[Dcache.scala 19:24]
  reg [3:0] offset_207; // @[Dcache.scala 19:24]
  reg [3:0] offset_208; // @[Dcache.scala 19:24]
  reg [3:0] offset_209; // @[Dcache.scala 19:24]
  reg [3:0] offset_210; // @[Dcache.scala 19:24]
  reg [3:0] offset_211; // @[Dcache.scala 19:24]
  reg [3:0] offset_212; // @[Dcache.scala 19:24]
  reg [3:0] offset_213; // @[Dcache.scala 19:24]
  reg [3:0] offset_214; // @[Dcache.scala 19:24]
  reg [3:0] offset_215; // @[Dcache.scala 19:24]
  reg [3:0] offset_216; // @[Dcache.scala 19:24]
  reg [3:0] offset_217; // @[Dcache.scala 19:24]
  reg [3:0] offset_218; // @[Dcache.scala 19:24]
  reg [3:0] offset_219; // @[Dcache.scala 19:24]
  reg [3:0] offset_220; // @[Dcache.scala 19:24]
  reg [3:0] offset_221; // @[Dcache.scala 19:24]
  reg [3:0] offset_222; // @[Dcache.scala 19:24]
  reg [3:0] offset_223; // @[Dcache.scala 19:24]
  reg [3:0] offset_224; // @[Dcache.scala 19:24]
  reg [3:0] offset_225; // @[Dcache.scala 19:24]
  reg [3:0] offset_226; // @[Dcache.scala 19:24]
  reg [3:0] offset_227; // @[Dcache.scala 19:24]
  reg [3:0] offset_228; // @[Dcache.scala 19:24]
  reg [3:0] offset_229; // @[Dcache.scala 19:24]
  reg [3:0] offset_230; // @[Dcache.scala 19:24]
  reg [3:0] offset_231; // @[Dcache.scala 19:24]
  reg [3:0] offset_232; // @[Dcache.scala 19:24]
  reg [3:0] offset_233; // @[Dcache.scala 19:24]
  reg [3:0] offset_234; // @[Dcache.scala 19:24]
  reg [3:0] offset_235; // @[Dcache.scala 19:24]
  reg [3:0] offset_236; // @[Dcache.scala 19:24]
  reg [3:0] offset_237; // @[Dcache.scala 19:24]
  reg [3:0] offset_238; // @[Dcache.scala 19:24]
  reg [3:0] offset_239; // @[Dcache.scala 19:24]
  reg [3:0] offset_240; // @[Dcache.scala 19:24]
  reg [3:0] offset_241; // @[Dcache.scala 19:24]
  reg [3:0] offset_242; // @[Dcache.scala 19:24]
  reg [3:0] offset_243; // @[Dcache.scala 19:24]
  reg [3:0] offset_244; // @[Dcache.scala 19:24]
  reg [3:0] offset_245; // @[Dcache.scala 19:24]
  reg [3:0] offset_246; // @[Dcache.scala 19:24]
  reg [3:0] offset_247; // @[Dcache.scala 19:24]
  reg [3:0] offset_248; // @[Dcache.scala 19:24]
  reg [3:0] offset_249; // @[Dcache.scala 19:24]
  reg [3:0] offset_250; // @[Dcache.scala 19:24]
  reg [3:0] offset_251; // @[Dcache.scala 19:24]
  reg [3:0] offset_252; // @[Dcache.scala 19:24]
  reg [3:0] offset_253; // @[Dcache.scala 19:24]
  reg [3:0] offset_254; // @[Dcache.scala 19:24]
  reg [3:0] offset_255; // @[Dcache.scala 19:24]
  reg [2:0] state; // @[Dcache.scala 26:22]
  wire [19:0] req_tag = io_dmem_data_addr[31:12]; // @[Dcache.scala 28:30]
  wire [7:0] req_index = io_dmem_data_addr[11:4]; // @[Dcache.scala 29:30]
  wire [3:0] req_offset = io_dmem_data_addr[3:0]; // @[Dcache.scala 30:30]
  wire [19:0] _GEN_1 = 8'h1 == req_index ? tag_1 : tag_0; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_2 = 8'h2 == req_index ? tag_2 : _GEN_1; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_3 = 8'h3 == req_index ? tag_3 : _GEN_2; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_4 = 8'h4 == req_index ? tag_4 : _GEN_3; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_5 = 8'h5 == req_index ? tag_5 : _GEN_4; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_6 = 8'h6 == req_index ? tag_6 : _GEN_5; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_7 = 8'h7 == req_index ? tag_7 : _GEN_6; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_8 = 8'h8 == req_index ? tag_8 : _GEN_7; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_9 = 8'h9 == req_index ? tag_9 : _GEN_8; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_10 = 8'ha == req_index ? tag_10 : _GEN_9; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_11 = 8'hb == req_index ? tag_11 : _GEN_10; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_12 = 8'hc == req_index ? tag_12 : _GEN_11; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_13 = 8'hd == req_index ? tag_13 : _GEN_12; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_14 = 8'he == req_index ? tag_14 : _GEN_13; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_15 = 8'hf == req_index ? tag_15 : _GEN_14; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_16 = 8'h10 == req_index ? tag_16 : _GEN_15; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_17 = 8'h11 == req_index ? tag_17 : _GEN_16; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_18 = 8'h12 == req_index ? tag_18 : _GEN_17; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_19 = 8'h13 == req_index ? tag_19 : _GEN_18; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_20 = 8'h14 == req_index ? tag_20 : _GEN_19; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_21 = 8'h15 == req_index ? tag_21 : _GEN_20; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_22 = 8'h16 == req_index ? tag_22 : _GEN_21; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_23 = 8'h17 == req_index ? tag_23 : _GEN_22; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_24 = 8'h18 == req_index ? tag_24 : _GEN_23; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_25 = 8'h19 == req_index ? tag_25 : _GEN_24; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_26 = 8'h1a == req_index ? tag_26 : _GEN_25; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_27 = 8'h1b == req_index ? tag_27 : _GEN_26; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_28 = 8'h1c == req_index ? tag_28 : _GEN_27; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_29 = 8'h1d == req_index ? tag_29 : _GEN_28; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_30 = 8'h1e == req_index ? tag_30 : _GEN_29; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_31 = 8'h1f == req_index ? tag_31 : _GEN_30; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_32 = 8'h20 == req_index ? tag_32 : _GEN_31; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_33 = 8'h21 == req_index ? tag_33 : _GEN_32; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_34 = 8'h22 == req_index ? tag_34 : _GEN_33; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_35 = 8'h23 == req_index ? tag_35 : _GEN_34; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_36 = 8'h24 == req_index ? tag_36 : _GEN_35; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_37 = 8'h25 == req_index ? tag_37 : _GEN_36; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_38 = 8'h26 == req_index ? tag_38 : _GEN_37; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_39 = 8'h27 == req_index ? tag_39 : _GEN_38; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_40 = 8'h28 == req_index ? tag_40 : _GEN_39; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_41 = 8'h29 == req_index ? tag_41 : _GEN_40; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_42 = 8'h2a == req_index ? tag_42 : _GEN_41; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_43 = 8'h2b == req_index ? tag_43 : _GEN_42; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_44 = 8'h2c == req_index ? tag_44 : _GEN_43; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_45 = 8'h2d == req_index ? tag_45 : _GEN_44; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_46 = 8'h2e == req_index ? tag_46 : _GEN_45; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_47 = 8'h2f == req_index ? tag_47 : _GEN_46; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_48 = 8'h30 == req_index ? tag_48 : _GEN_47; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_49 = 8'h31 == req_index ? tag_49 : _GEN_48; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_50 = 8'h32 == req_index ? tag_50 : _GEN_49; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_51 = 8'h33 == req_index ? tag_51 : _GEN_50; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_52 = 8'h34 == req_index ? tag_52 : _GEN_51; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_53 = 8'h35 == req_index ? tag_53 : _GEN_52; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_54 = 8'h36 == req_index ? tag_54 : _GEN_53; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_55 = 8'h37 == req_index ? tag_55 : _GEN_54; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_56 = 8'h38 == req_index ? tag_56 : _GEN_55; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_57 = 8'h39 == req_index ? tag_57 : _GEN_56; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_58 = 8'h3a == req_index ? tag_58 : _GEN_57; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_59 = 8'h3b == req_index ? tag_59 : _GEN_58; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_60 = 8'h3c == req_index ? tag_60 : _GEN_59; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_61 = 8'h3d == req_index ? tag_61 : _GEN_60; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_62 = 8'h3e == req_index ? tag_62 : _GEN_61; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_63 = 8'h3f == req_index ? tag_63 : _GEN_62; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_64 = 8'h40 == req_index ? tag_64 : _GEN_63; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_65 = 8'h41 == req_index ? tag_65 : _GEN_64; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_66 = 8'h42 == req_index ? tag_66 : _GEN_65; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_67 = 8'h43 == req_index ? tag_67 : _GEN_66; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_68 = 8'h44 == req_index ? tag_68 : _GEN_67; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_69 = 8'h45 == req_index ? tag_69 : _GEN_68; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_70 = 8'h46 == req_index ? tag_70 : _GEN_69; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_71 = 8'h47 == req_index ? tag_71 : _GEN_70; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_72 = 8'h48 == req_index ? tag_72 : _GEN_71; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_73 = 8'h49 == req_index ? tag_73 : _GEN_72; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_74 = 8'h4a == req_index ? tag_74 : _GEN_73; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_75 = 8'h4b == req_index ? tag_75 : _GEN_74; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_76 = 8'h4c == req_index ? tag_76 : _GEN_75; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_77 = 8'h4d == req_index ? tag_77 : _GEN_76; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_78 = 8'h4e == req_index ? tag_78 : _GEN_77; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_79 = 8'h4f == req_index ? tag_79 : _GEN_78; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_80 = 8'h50 == req_index ? tag_80 : _GEN_79; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_81 = 8'h51 == req_index ? tag_81 : _GEN_80; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_82 = 8'h52 == req_index ? tag_82 : _GEN_81; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_83 = 8'h53 == req_index ? tag_83 : _GEN_82; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_84 = 8'h54 == req_index ? tag_84 : _GEN_83; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_85 = 8'h55 == req_index ? tag_85 : _GEN_84; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_86 = 8'h56 == req_index ? tag_86 : _GEN_85; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_87 = 8'h57 == req_index ? tag_87 : _GEN_86; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_88 = 8'h58 == req_index ? tag_88 : _GEN_87; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_89 = 8'h59 == req_index ? tag_89 : _GEN_88; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_90 = 8'h5a == req_index ? tag_90 : _GEN_89; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_91 = 8'h5b == req_index ? tag_91 : _GEN_90; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_92 = 8'h5c == req_index ? tag_92 : _GEN_91; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_93 = 8'h5d == req_index ? tag_93 : _GEN_92; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_94 = 8'h5e == req_index ? tag_94 : _GEN_93; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_95 = 8'h5f == req_index ? tag_95 : _GEN_94; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_96 = 8'h60 == req_index ? tag_96 : _GEN_95; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_97 = 8'h61 == req_index ? tag_97 : _GEN_96; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_98 = 8'h62 == req_index ? tag_98 : _GEN_97; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_99 = 8'h63 == req_index ? tag_99 : _GEN_98; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_100 = 8'h64 == req_index ? tag_100 : _GEN_99; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_101 = 8'h65 == req_index ? tag_101 : _GEN_100; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_102 = 8'h66 == req_index ? tag_102 : _GEN_101; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_103 = 8'h67 == req_index ? tag_103 : _GEN_102; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_104 = 8'h68 == req_index ? tag_104 : _GEN_103; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_105 = 8'h69 == req_index ? tag_105 : _GEN_104; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_106 = 8'h6a == req_index ? tag_106 : _GEN_105; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_107 = 8'h6b == req_index ? tag_107 : _GEN_106; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_108 = 8'h6c == req_index ? tag_108 : _GEN_107; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_109 = 8'h6d == req_index ? tag_109 : _GEN_108; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_110 = 8'h6e == req_index ? tag_110 : _GEN_109; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_111 = 8'h6f == req_index ? tag_111 : _GEN_110; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_112 = 8'h70 == req_index ? tag_112 : _GEN_111; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_113 = 8'h71 == req_index ? tag_113 : _GEN_112; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_114 = 8'h72 == req_index ? tag_114 : _GEN_113; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_115 = 8'h73 == req_index ? tag_115 : _GEN_114; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_116 = 8'h74 == req_index ? tag_116 : _GEN_115; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_117 = 8'h75 == req_index ? tag_117 : _GEN_116; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_118 = 8'h76 == req_index ? tag_118 : _GEN_117; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_119 = 8'h77 == req_index ? tag_119 : _GEN_118; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_120 = 8'h78 == req_index ? tag_120 : _GEN_119; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_121 = 8'h79 == req_index ? tag_121 : _GEN_120; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_122 = 8'h7a == req_index ? tag_122 : _GEN_121; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_123 = 8'h7b == req_index ? tag_123 : _GEN_122; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_124 = 8'h7c == req_index ? tag_124 : _GEN_123; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_125 = 8'h7d == req_index ? tag_125 : _GEN_124; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_126 = 8'h7e == req_index ? tag_126 : _GEN_125; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_127 = 8'h7f == req_index ? tag_127 : _GEN_126; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_128 = 8'h80 == req_index ? tag_128 : _GEN_127; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_129 = 8'h81 == req_index ? tag_129 : _GEN_128; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_130 = 8'h82 == req_index ? tag_130 : _GEN_129; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_131 = 8'h83 == req_index ? tag_131 : _GEN_130; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_132 = 8'h84 == req_index ? tag_132 : _GEN_131; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_133 = 8'h85 == req_index ? tag_133 : _GEN_132; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_134 = 8'h86 == req_index ? tag_134 : _GEN_133; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_135 = 8'h87 == req_index ? tag_135 : _GEN_134; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_136 = 8'h88 == req_index ? tag_136 : _GEN_135; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_137 = 8'h89 == req_index ? tag_137 : _GEN_136; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_138 = 8'h8a == req_index ? tag_138 : _GEN_137; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_139 = 8'h8b == req_index ? tag_139 : _GEN_138; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_140 = 8'h8c == req_index ? tag_140 : _GEN_139; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_141 = 8'h8d == req_index ? tag_141 : _GEN_140; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_142 = 8'h8e == req_index ? tag_142 : _GEN_141; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_143 = 8'h8f == req_index ? tag_143 : _GEN_142; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_144 = 8'h90 == req_index ? tag_144 : _GEN_143; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_145 = 8'h91 == req_index ? tag_145 : _GEN_144; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_146 = 8'h92 == req_index ? tag_146 : _GEN_145; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_147 = 8'h93 == req_index ? tag_147 : _GEN_146; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_148 = 8'h94 == req_index ? tag_148 : _GEN_147; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_149 = 8'h95 == req_index ? tag_149 : _GEN_148; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_150 = 8'h96 == req_index ? tag_150 : _GEN_149; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_151 = 8'h97 == req_index ? tag_151 : _GEN_150; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_152 = 8'h98 == req_index ? tag_152 : _GEN_151; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_153 = 8'h99 == req_index ? tag_153 : _GEN_152; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_154 = 8'h9a == req_index ? tag_154 : _GEN_153; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_155 = 8'h9b == req_index ? tag_155 : _GEN_154; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_156 = 8'h9c == req_index ? tag_156 : _GEN_155; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_157 = 8'h9d == req_index ? tag_157 : _GEN_156; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_158 = 8'h9e == req_index ? tag_158 : _GEN_157; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_159 = 8'h9f == req_index ? tag_159 : _GEN_158; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_160 = 8'ha0 == req_index ? tag_160 : _GEN_159; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_161 = 8'ha1 == req_index ? tag_161 : _GEN_160; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_162 = 8'ha2 == req_index ? tag_162 : _GEN_161; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_163 = 8'ha3 == req_index ? tag_163 : _GEN_162; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_164 = 8'ha4 == req_index ? tag_164 : _GEN_163; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_165 = 8'ha5 == req_index ? tag_165 : _GEN_164; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_166 = 8'ha6 == req_index ? tag_166 : _GEN_165; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_167 = 8'ha7 == req_index ? tag_167 : _GEN_166; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_168 = 8'ha8 == req_index ? tag_168 : _GEN_167; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_169 = 8'ha9 == req_index ? tag_169 : _GEN_168; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_170 = 8'haa == req_index ? tag_170 : _GEN_169; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_171 = 8'hab == req_index ? tag_171 : _GEN_170; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_172 = 8'hac == req_index ? tag_172 : _GEN_171; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_173 = 8'had == req_index ? tag_173 : _GEN_172; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_174 = 8'hae == req_index ? tag_174 : _GEN_173; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_175 = 8'haf == req_index ? tag_175 : _GEN_174; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_176 = 8'hb0 == req_index ? tag_176 : _GEN_175; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_177 = 8'hb1 == req_index ? tag_177 : _GEN_176; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_178 = 8'hb2 == req_index ? tag_178 : _GEN_177; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_179 = 8'hb3 == req_index ? tag_179 : _GEN_178; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_180 = 8'hb4 == req_index ? tag_180 : _GEN_179; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_181 = 8'hb5 == req_index ? tag_181 : _GEN_180; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_182 = 8'hb6 == req_index ? tag_182 : _GEN_181; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_183 = 8'hb7 == req_index ? tag_183 : _GEN_182; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_184 = 8'hb8 == req_index ? tag_184 : _GEN_183; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_185 = 8'hb9 == req_index ? tag_185 : _GEN_184; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_186 = 8'hba == req_index ? tag_186 : _GEN_185; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_187 = 8'hbb == req_index ? tag_187 : _GEN_186; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_188 = 8'hbc == req_index ? tag_188 : _GEN_187; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_189 = 8'hbd == req_index ? tag_189 : _GEN_188; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_190 = 8'hbe == req_index ? tag_190 : _GEN_189; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_191 = 8'hbf == req_index ? tag_191 : _GEN_190; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_192 = 8'hc0 == req_index ? tag_192 : _GEN_191; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_193 = 8'hc1 == req_index ? tag_193 : _GEN_192; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_194 = 8'hc2 == req_index ? tag_194 : _GEN_193; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_195 = 8'hc3 == req_index ? tag_195 : _GEN_194; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_196 = 8'hc4 == req_index ? tag_196 : _GEN_195; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_197 = 8'hc5 == req_index ? tag_197 : _GEN_196; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_198 = 8'hc6 == req_index ? tag_198 : _GEN_197; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_199 = 8'hc7 == req_index ? tag_199 : _GEN_198; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_200 = 8'hc8 == req_index ? tag_200 : _GEN_199; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_201 = 8'hc9 == req_index ? tag_201 : _GEN_200; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_202 = 8'hca == req_index ? tag_202 : _GEN_201; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_203 = 8'hcb == req_index ? tag_203 : _GEN_202; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_204 = 8'hcc == req_index ? tag_204 : _GEN_203; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_205 = 8'hcd == req_index ? tag_205 : _GEN_204; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_206 = 8'hce == req_index ? tag_206 : _GEN_205; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_207 = 8'hcf == req_index ? tag_207 : _GEN_206; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_208 = 8'hd0 == req_index ? tag_208 : _GEN_207; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_209 = 8'hd1 == req_index ? tag_209 : _GEN_208; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_210 = 8'hd2 == req_index ? tag_210 : _GEN_209; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_211 = 8'hd3 == req_index ? tag_211 : _GEN_210; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_212 = 8'hd4 == req_index ? tag_212 : _GEN_211; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_213 = 8'hd5 == req_index ? tag_213 : _GEN_212; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_214 = 8'hd6 == req_index ? tag_214 : _GEN_213; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_215 = 8'hd7 == req_index ? tag_215 : _GEN_214; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_216 = 8'hd8 == req_index ? tag_216 : _GEN_215; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_217 = 8'hd9 == req_index ? tag_217 : _GEN_216; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_218 = 8'hda == req_index ? tag_218 : _GEN_217; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_219 = 8'hdb == req_index ? tag_219 : _GEN_218; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_220 = 8'hdc == req_index ? tag_220 : _GEN_219; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_221 = 8'hdd == req_index ? tag_221 : _GEN_220; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_222 = 8'hde == req_index ? tag_222 : _GEN_221; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_223 = 8'hdf == req_index ? tag_223 : _GEN_222; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_224 = 8'he0 == req_index ? tag_224 : _GEN_223; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_225 = 8'he1 == req_index ? tag_225 : _GEN_224; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_226 = 8'he2 == req_index ? tag_226 : _GEN_225; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_227 = 8'he3 == req_index ? tag_227 : _GEN_226; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_228 = 8'he4 == req_index ? tag_228 : _GEN_227; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_229 = 8'he5 == req_index ? tag_229 : _GEN_228; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_230 = 8'he6 == req_index ? tag_230 : _GEN_229; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_231 = 8'he7 == req_index ? tag_231 : _GEN_230; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_232 = 8'he8 == req_index ? tag_232 : _GEN_231; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_233 = 8'he9 == req_index ? tag_233 : _GEN_232; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_234 = 8'hea == req_index ? tag_234 : _GEN_233; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_235 = 8'heb == req_index ? tag_235 : _GEN_234; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_236 = 8'hec == req_index ? tag_236 : _GEN_235; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_237 = 8'hed == req_index ? tag_237 : _GEN_236; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_238 = 8'hee == req_index ? tag_238 : _GEN_237; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_239 = 8'hef == req_index ? tag_239 : _GEN_238; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_240 = 8'hf0 == req_index ? tag_240 : _GEN_239; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_241 = 8'hf1 == req_index ? tag_241 : _GEN_240; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_242 = 8'hf2 == req_index ? tag_242 : _GEN_241; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_243 = 8'hf3 == req_index ? tag_243 : _GEN_242; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_244 = 8'hf4 == req_index ? tag_244 : _GEN_243; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_245 = 8'hf5 == req_index ? tag_245 : _GEN_244; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_246 = 8'hf6 == req_index ? tag_246 : _GEN_245; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_247 = 8'hf7 == req_index ? tag_247 : _GEN_246; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_248 = 8'hf8 == req_index ? tag_248 : _GEN_247; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_249 = 8'hf9 == req_index ? tag_249 : _GEN_248; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_250 = 8'hfa == req_index ? tag_250 : _GEN_249; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_251 = 8'hfb == req_index ? tag_251 : _GEN_250; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_252 = 8'hfc == req_index ? tag_252 : _GEN_251; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_253 = 8'hfd == req_index ? tag_253 : _GEN_252; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_254 = 8'hfe == req_index ? tag_254 : _GEN_253; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire [19:0] _GEN_255 = 8'hff == req_index ? tag_255 : _GEN_254; // @[Dcache.scala 34:36 Dcache.scala 34:36]
  wire  _GEN_257 = 8'h1 == req_index ? valid_1 : valid_0; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_258 = 8'h2 == req_index ? valid_2 : _GEN_257; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_259 = 8'h3 == req_index ? valid_3 : _GEN_258; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_260 = 8'h4 == req_index ? valid_4 : _GEN_259; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_261 = 8'h5 == req_index ? valid_5 : _GEN_260; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_262 = 8'h6 == req_index ? valid_6 : _GEN_261; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_263 = 8'h7 == req_index ? valid_7 : _GEN_262; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_264 = 8'h8 == req_index ? valid_8 : _GEN_263; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_265 = 8'h9 == req_index ? valid_9 : _GEN_264; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_266 = 8'ha == req_index ? valid_10 : _GEN_265; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_267 = 8'hb == req_index ? valid_11 : _GEN_266; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_268 = 8'hc == req_index ? valid_12 : _GEN_267; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_269 = 8'hd == req_index ? valid_13 : _GEN_268; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_270 = 8'he == req_index ? valid_14 : _GEN_269; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_271 = 8'hf == req_index ? valid_15 : _GEN_270; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_272 = 8'h10 == req_index ? valid_16 : _GEN_271; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_273 = 8'h11 == req_index ? valid_17 : _GEN_272; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_274 = 8'h12 == req_index ? valid_18 : _GEN_273; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_275 = 8'h13 == req_index ? valid_19 : _GEN_274; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_276 = 8'h14 == req_index ? valid_20 : _GEN_275; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_277 = 8'h15 == req_index ? valid_21 : _GEN_276; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_278 = 8'h16 == req_index ? valid_22 : _GEN_277; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_279 = 8'h17 == req_index ? valid_23 : _GEN_278; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_280 = 8'h18 == req_index ? valid_24 : _GEN_279; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_281 = 8'h19 == req_index ? valid_25 : _GEN_280; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_282 = 8'h1a == req_index ? valid_26 : _GEN_281; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_283 = 8'h1b == req_index ? valid_27 : _GEN_282; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_284 = 8'h1c == req_index ? valid_28 : _GEN_283; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_285 = 8'h1d == req_index ? valid_29 : _GEN_284; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_286 = 8'h1e == req_index ? valid_30 : _GEN_285; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_287 = 8'h1f == req_index ? valid_31 : _GEN_286; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_288 = 8'h20 == req_index ? valid_32 : _GEN_287; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_289 = 8'h21 == req_index ? valid_33 : _GEN_288; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_290 = 8'h22 == req_index ? valid_34 : _GEN_289; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_291 = 8'h23 == req_index ? valid_35 : _GEN_290; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_292 = 8'h24 == req_index ? valid_36 : _GEN_291; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_293 = 8'h25 == req_index ? valid_37 : _GEN_292; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_294 = 8'h26 == req_index ? valid_38 : _GEN_293; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_295 = 8'h27 == req_index ? valid_39 : _GEN_294; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_296 = 8'h28 == req_index ? valid_40 : _GEN_295; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_297 = 8'h29 == req_index ? valid_41 : _GEN_296; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_298 = 8'h2a == req_index ? valid_42 : _GEN_297; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_299 = 8'h2b == req_index ? valid_43 : _GEN_298; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_300 = 8'h2c == req_index ? valid_44 : _GEN_299; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_301 = 8'h2d == req_index ? valid_45 : _GEN_300; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_302 = 8'h2e == req_index ? valid_46 : _GEN_301; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_303 = 8'h2f == req_index ? valid_47 : _GEN_302; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_304 = 8'h30 == req_index ? valid_48 : _GEN_303; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_305 = 8'h31 == req_index ? valid_49 : _GEN_304; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_306 = 8'h32 == req_index ? valid_50 : _GEN_305; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_307 = 8'h33 == req_index ? valid_51 : _GEN_306; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_308 = 8'h34 == req_index ? valid_52 : _GEN_307; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_309 = 8'h35 == req_index ? valid_53 : _GEN_308; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_310 = 8'h36 == req_index ? valid_54 : _GEN_309; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_311 = 8'h37 == req_index ? valid_55 : _GEN_310; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_312 = 8'h38 == req_index ? valid_56 : _GEN_311; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_313 = 8'h39 == req_index ? valid_57 : _GEN_312; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_314 = 8'h3a == req_index ? valid_58 : _GEN_313; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_315 = 8'h3b == req_index ? valid_59 : _GEN_314; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_316 = 8'h3c == req_index ? valid_60 : _GEN_315; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_317 = 8'h3d == req_index ? valid_61 : _GEN_316; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_318 = 8'h3e == req_index ? valid_62 : _GEN_317; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_319 = 8'h3f == req_index ? valid_63 : _GEN_318; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_320 = 8'h40 == req_index ? valid_64 : _GEN_319; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_321 = 8'h41 == req_index ? valid_65 : _GEN_320; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_322 = 8'h42 == req_index ? valid_66 : _GEN_321; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_323 = 8'h43 == req_index ? valid_67 : _GEN_322; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_324 = 8'h44 == req_index ? valid_68 : _GEN_323; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_325 = 8'h45 == req_index ? valid_69 : _GEN_324; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_326 = 8'h46 == req_index ? valid_70 : _GEN_325; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_327 = 8'h47 == req_index ? valid_71 : _GEN_326; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_328 = 8'h48 == req_index ? valid_72 : _GEN_327; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_329 = 8'h49 == req_index ? valid_73 : _GEN_328; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_330 = 8'h4a == req_index ? valid_74 : _GEN_329; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_331 = 8'h4b == req_index ? valid_75 : _GEN_330; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_332 = 8'h4c == req_index ? valid_76 : _GEN_331; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_333 = 8'h4d == req_index ? valid_77 : _GEN_332; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_334 = 8'h4e == req_index ? valid_78 : _GEN_333; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_335 = 8'h4f == req_index ? valid_79 : _GEN_334; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_336 = 8'h50 == req_index ? valid_80 : _GEN_335; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_337 = 8'h51 == req_index ? valid_81 : _GEN_336; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_338 = 8'h52 == req_index ? valid_82 : _GEN_337; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_339 = 8'h53 == req_index ? valid_83 : _GEN_338; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_340 = 8'h54 == req_index ? valid_84 : _GEN_339; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_341 = 8'h55 == req_index ? valid_85 : _GEN_340; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_342 = 8'h56 == req_index ? valid_86 : _GEN_341; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_343 = 8'h57 == req_index ? valid_87 : _GEN_342; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_344 = 8'h58 == req_index ? valid_88 : _GEN_343; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_345 = 8'h59 == req_index ? valid_89 : _GEN_344; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_346 = 8'h5a == req_index ? valid_90 : _GEN_345; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_347 = 8'h5b == req_index ? valid_91 : _GEN_346; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_348 = 8'h5c == req_index ? valid_92 : _GEN_347; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_349 = 8'h5d == req_index ? valid_93 : _GEN_348; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_350 = 8'h5e == req_index ? valid_94 : _GEN_349; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_351 = 8'h5f == req_index ? valid_95 : _GEN_350; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_352 = 8'h60 == req_index ? valid_96 : _GEN_351; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_353 = 8'h61 == req_index ? valid_97 : _GEN_352; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_354 = 8'h62 == req_index ? valid_98 : _GEN_353; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_355 = 8'h63 == req_index ? valid_99 : _GEN_354; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_356 = 8'h64 == req_index ? valid_100 : _GEN_355; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_357 = 8'h65 == req_index ? valid_101 : _GEN_356; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_358 = 8'h66 == req_index ? valid_102 : _GEN_357; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_359 = 8'h67 == req_index ? valid_103 : _GEN_358; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_360 = 8'h68 == req_index ? valid_104 : _GEN_359; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_361 = 8'h69 == req_index ? valid_105 : _GEN_360; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_362 = 8'h6a == req_index ? valid_106 : _GEN_361; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_363 = 8'h6b == req_index ? valid_107 : _GEN_362; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_364 = 8'h6c == req_index ? valid_108 : _GEN_363; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_365 = 8'h6d == req_index ? valid_109 : _GEN_364; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_366 = 8'h6e == req_index ? valid_110 : _GEN_365; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_367 = 8'h6f == req_index ? valid_111 : _GEN_366; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_368 = 8'h70 == req_index ? valid_112 : _GEN_367; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_369 = 8'h71 == req_index ? valid_113 : _GEN_368; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_370 = 8'h72 == req_index ? valid_114 : _GEN_369; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_371 = 8'h73 == req_index ? valid_115 : _GEN_370; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_372 = 8'h74 == req_index ? valid_116 : _GEN_371; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_373 = 8'h75 == req_index ? valid_117 : _GEN_372; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_374 = 8'h76 == req_index ? valid_118 : _GEN_373; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_375 = 8'h77 == req_index ? valid_119 : _GEN_374; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_376 = 8'h78 == req_index ? valid_120 : _GEN_375; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_377 = 8'h79 == req_index ? valid_121 : _GEN_376; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_378 = 8'h7a == req_index ? valid_122 : _GEN_377; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_379 = 8'h7b == req_index ? valid_123 : _GEN_378; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_380 = 8'h7c == req_index ? valid_124 : _GEN_379; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_381 = 8'h7d == req_index ? valid_125 : _GEN_380; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_382 = 8'h7e == req_index ? valid_126 : _GEN_381; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_383 = 8'h7f == req_index ? valid_127 : _GEN_382; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_384 = 8'h80 == req_index ? valid_128 : _GEN_383; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_385 = 8'h81 == req_index ? valid_129 : _GEN_384; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_386 = 8'h82 == req_index ? valid_130 : _GEN_385; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_387 = 8'h83 == req_index ? valid_131 : _GEN_386; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_388 = 8'h84 == req_index ? valid_132 : _GEN_387; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_389 = 8'h85 == req_index ? valid_133 : _GEN_388; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_390 = 8'h86 == req_index ? valid_134 : _GEN_389; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_391 = 8'h87 == req_index ? valid_135 : _GEN_390; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_392 = 8'h88 == req_index ? valid_136 : _GEN_391; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_393 = 8'h89 == req_index ? valid_137 : _GEN_392; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_394 = 8'h8a == req_index ? valid_138 : _GEN_393; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_395 = 8'h8b == req_index ? valid_139 : _GEN_394; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_396 = 8'h8c == req_index ? valid_140 : _GEN_395; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_397 = 8'h8d == req_index ? valid_141 : _GEN_396; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_398 = 8'h8e == req_index ? valid_142 : _GEN_397; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_399 = 8'h8f == req_index ? valid_143 : _GEN_398; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_400 = 8'h90 == req_index ? valid_144 : _GEN_399; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_401 = 8'h91 == req_index ? valid_145 : _GEN_400; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_402 = 8'h92 == req_index ? valid_146 : _GEN_401; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_403 = 8'h93 == req_index ? valid_147 : _GEN_402; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_404 = 8'h94 == req_index ? valid_148 : _GEN_403; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_405 = 8'h95 == req_index ? valid_149 : _GEN_404; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_406 = 8'h96 == req_index ? valid_150 : _GEN_405; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_407 = 8'h97 == req_index ? valid_151 : _GEN_406; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_408 = 8'h98 == req_index ? valid_152 : _GEN_407; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_409 = 8'h99 == req_index ? valid_153 : _GEN_408; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_410 = 8'h9a == req_index ? valid_154 : _GEN_409; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_411 = 8'h9b == req_index ? valid_155 : _GEN_410; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_412 = 8'h9c == req_index ? valid_156 : _GEN_411; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_413 = 8'h9d == req_index ? valid_157 : _GEN_412; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_414 = 8'h9e == req_index ? valid_158 : _GEN_413; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_415 = 8'h9f == req_index ? valid_159 : _GEN_414; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_416 = 8'ha0 == req_index ? valid_160 : _GEN_415; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_417 = 8'ha1 == req_index ? valid_161 : _GEN_416; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_418 = 8'ha2 == req_index ? valid_162 : _GEN_417; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_419 = 8'ha3 == req_index ? valid_163 : _GEN_418; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_420 = 8'ha4 == req_index ? valid_164 : _GEN_419; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_421 = 8'ha5 == req_index ? valid_165 : _GEN_420; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_422 = 8'ha6 == req_index ? valid_166 : _GEN_421; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_423 = 8'ha7 == req_index ? valid_167 : _GEN_422; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_424 = 8'ha8 == req_index ? valid_168 : _GEN_423; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_425 = 8'ha9 == req_index ? valid_169 : _GEN_424; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_426 = 8'haa == req_index ? valid_170 : _GEN_425; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_427 = 8'hab == req_index ? valid_171 : _GEN_426; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_428 = 8'hac == req_index ? valid_172 : _GEN_427; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_429 = 8'had == req_index ? valid_173 : _GEN_428; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_430 = 8'hae == req_index ? valid_174 : _GEN_429; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_431 = 8'haf == req_index ? valid_175 : _GEN_430; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_432 = 8'hb0 == req_index ? valid_176 : _GEN_431; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_433 = 8'hb1 == req_index ? valid_177 : _GEN_432; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_434 = 8'hb2 == req_index ? valid_178 : _GEN_433; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_435 = 8'hb3 == req_index ? valid_179 : _GEN_434; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_436 = 8'hb4 == req_index ? valid_180 : _GEN_435; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_437 = 8'hb5 == req_index ? valid_181 : _GEN_436; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_438 = 8'hb6 == req_index ? valid_182 : _GEN_437; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_439 = 8'hb7 == req_index ? valid_183 : _GEN_438; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_440 = 8'hb8 == req_index ? valid_184 : _GEN_439; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_441 = 8'hb9 == req_index ? valid_185 : _GEN_440; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_442 = 8'hba == req_index ? valid_186 : _GEN_441; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_443 = 8'hbb == req_index ? valid_187 : _GEN_442; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_444 = 8'hbc == req_index ? valid_188 : _GEN_443; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_445 = 8'hbd == req_index ? valid_189 : _GEN_444; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_446 = 8'hbe == req_index ? valid_190 : _GEN_445; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_447 = 8'hbf == req_index ? valid_191 : _GEN_446; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_448 = 8'hc0 == req_index ? valid_192 : _GEN_447; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_449 = 8'hc1 == req_index ? valid_193 : _GEN_448; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_450 = 8'hc2 == req_index ? valid_194 : _GEN_449; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_451 = 8'hc3 == req_index ? valid_195 : _GEN_450; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_452 = 8'hc4 == req_index ? valid_196 : _GEN_451; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_453 = 8'hc5 == req_index ? valid_197 : _GEN_452; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_454 = 8'hc6 == req_index ? valid_198 : _GEN_453; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_455 = 8'hc7 == req_index ? valid_199 : _GEN_454; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_456 = 8'hc8 == req_index ? valid_200 : _GEN_455; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_457 = 8'hc9 == req_index ? valid_201 : _GEN_456; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_458 = 8'hca == req_index ? valid_202 : _GEN_457; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_459 = 8'hcb == req_index ? valid_203 : _GEN_458; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_460 = 8'hcc == req_index ? valid_204 : _GEN_459; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_461 = 8'hcd == req_index ? valid_205 : _GEN_460; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_462 = 8'hce == req_index ? valid_206 : _GEN_461; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_463 = 8'hcf == req_index ? valid_207 : _GEN_462; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_464 = 8'hd0 == req_index ? valid_208 : _GEN_463; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_465 = 8'hd1 == req_index ? valid_209 : _GEN_464; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_466 = 8'hd2 == req_index ? valid_210 : _GEN_465; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_467 = 8'hd3 == req_index ? valid_211 : _GEN_466; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_468 = 8'hd4 == req_index ? valid_212 : _GEN_467; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_469 = 8'hd5 == req_index ? valid_213 : _GEN_468; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_470 = 8'hd6 == req_index ? valid_214 : _GEN_469; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_471 = 8'hd7 == req_index ? valid_215 : _GEN_470; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_472 = 8'hd8 == req_index ? valid_216 : _GEN_471; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_473 = 8'hd9 == req_index ? valid_217 : _GEN_472; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_474 = 8'hda == req_index ? valid_218 : _GEN_473; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_475 = 8'hdb == req_index ? valid_219 : _GEN_474; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_476 = 8'hdc == req_index ? valid_220 : _GEN_475; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_477 = 8'hdd == req_index ? valid_221 : _GEN_476; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_478 = 8'hde == req_index ? valid_222 : _GEN_477; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_479 = 8'hdf == req_index ? valid_223 : _GEN_478; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_480 = 8'he0 == req_index ? valid_224 : _GEN_479; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_481 = 8'he1 == req_index ? valid_225 : _GEN_480; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_482 = 8'he2 == req_index ? valid_226 : _GEN_481; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_483 = 8'he3 == req_index ? valid_227 : _GEN_482; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_484 = 8'he4 == req_index ? valid_228 : _GEN_483; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_485 = 8'he5 == req_index ? valid_229 : _GEN_484; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_486 = 8'he6 == req_index ? valid_230 : _GEN_485; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_487 = 8'he7 == req_index ? valid_231 : _GEN_486; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_488 = 8'he8 == req_index ? valid_232 : _GEN_487; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_489 = 8'he9 == req_index ? valid_233 : _GEN_488; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_490 = 8'hea == req_index ? valid_234 : _GEN_489; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_491 = 8'heb == req_index ? valid_235 : _GEN_490; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_492 = 8'hec == req_index ? valid_236 : _GEN_491; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_493 = 8'hed == req_index ? valid_237 : _GEN_492; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_494 = 8'hee == req_index ? valid_238 : _GEN_493; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_495 = 8'hef == req_index ? valid_239 : _GEN_494; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_496 = 8'hf0 == req_index ? valid_240 : _GEN_495; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_497 = 8'hf1 == req_index ? valid_241 : _GEN_496; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_498 = 8'hf2 == req_index ? valid_242 : _GEN_497; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_499 = 8'hf3 == req_index ? valid_243 : _GEN_498; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_500 = 8'hf4 == req_index ? valid_244 : _GEN_499; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_501 = 8'hf5 == req_index ? valid_245 : _GEN_500; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_502 = 8'hf6 == req_index ? valid_246 : _GEN_501; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_503 = 8'hf7 == req_index ? valid_247 : _GEN_502; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_504 = 8'hf8 == req_index ? valid_248 : _GEN_503; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_505 = 8'hf9 == req_index ? valid_249 : _GEN_504; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_506 = 8'hfa == req_index ? valid_250 : _GEN_505; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_507 = 8'hfb == req_index ? valid_251 : _GEN_506; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_508 = 8'hfc == req_index ? valid_252 : _GEN_507; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_509 = 8'hfd == req_index ? valid_253 : _GEN_508; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_510 = 8'hfe == req_index ? valid_254 : _GEN_509; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _GEN_511 = 8'hff == req_index ? valid_255 : _GEN_510; // @[Dcache.scala 34:49 Dcache.scala 34:49]
  wire  _cache_hit_T_2 = state == 3'h1; // @[Dcache.scala 34:78]
  wire  cache_hit = _GEN_255 == req_tag & _GEN_511 & state == 3'h1; // @[Dcache.scala 34:69]
  wire  _GEN_513 = 8'h1 == req_index ? dirty_1 : dirty_0; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_514 = 8'h2 == req_index ? dirty_2 : _GEN_513; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_515 = 8'h3 == req_index ? dirty_3 : _GEN_514; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_516 = 8'h4 == req_index ? dirty_4 : _GEN_515; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_517 = 8'h5 == req_index ? dirty_5 : _GEN_516; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_518 = 8'h6 == req_index ? dirty_6 : _GEN_517; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_519 = 8'h7 == req_index ? dirty_7 : _GEN_518; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_520 = 8'h8 == req_index ? dirty_8 : _GEN_519; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_521 = 8'h9 == req_index ? dirty_9 : _GEN_520; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_522 = 8'ha == req_index ? dirty_10 : _GEN_521; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_523 = 8'hb == req_index ? dirty_11 : _GEN_522; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_524 = 8'hc == req_index ? dirty_12 : _GEN_523; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_525 = 8'hd == req_index ? dirty_13 : _GEN_524; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_526 = 8'he == req_index ? dirty_14 : _GEN_525; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_527 = 8'hf == req_index ? dirty_15 : _GEN_526; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_528 = 8'h10 == req_index ? dirty_16 : _GEN_527; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_529 = 8'h11 == req_index ? dirty_17 : _GEN_528; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_530 = 8'h12 == req_index ? dirty_18 : _GEN_529; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_531 = 8'h13 == req_index ? dirty_19 : _GEN_530; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_532 = 8'h14 == req_index ? dirty_20 : _GEN_531; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_533 = 8'h15 == req_index ? dirty_21 : _GEN_532; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_534 = 8'h16 == req_index ? dirty_22 : _GEN_533; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_535 = 8'h17 == req_index ? dirty_23 : _GEN_534; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_536 = 8'h18 == req_index ? dirty_24 : _GEN_535; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_537 = 8'h19 == req_index ? dirty_25 : _GEN_536; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_538 = 8'h1a == req_index ? dirty_26 : _GEN_537; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_539 = 8'h1b == req_index ? dirty_27 : _GEN_538; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_540 = 8'h1c == req_index ? dirty_28 : _GEN_539; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_541 = 8'h1d == req_index ? dirty_29 : _GEN_540; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_542 = 8'h1e == req_index ? dirty_30 : _GEN_541; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_543 = 8'h1f == req_index ? dirty_31 : _GEN_542; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_544 = 8'h20 == req_index ? dirty_32 : _GEN_543; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_545 = 8'h21 == req_index ? dirty_33 : _GEN_544; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_546 = 8'h22 == req_index ? dirty_34 : _GEN_545; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_547 = 8'h23 == req_index ? dirty_35 : _GEN_546; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_548 = 8'h24 == req_index ? dirty_36 : _GEN_547; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_549 = 8'h25 == req_index ? dirty_37 : _GEN_548; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_550 = 8'h26 == req_index ? dirty_38 : _GEN_549; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_551 = 8'h27 == req_index ? dirty_39 : _GEN_550; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_552 = 8'h28 == req_index ? dirty_40 : _GEN_551; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_553 = 8'h29 == req_index ? dirty_41 : _GEN_552; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_554 = 8'h2a == req_index ? dirty_42 : _GEN_553; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_555 = 8'h2b == req_index ? dirty_43 : _GEN_554; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_556 = 8'h2c == req_index ? dirty_44 : _GEN_555; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_557 = 8'h2d == req_index ? dirty_45 : _GEN_556; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_558 = 8'h2e == req_index ? dirty_46 : _GEN_557; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_559 = 8'h2f == req_index ? dirty_47 : _GEN_558; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_560 = 8'h30 == req_index ? dirty_48 : _GEN_559; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_561 = 8'h31 == req_index ? dirty_49 : _GEN_560; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_562 = 8'h32 == req_index ? dirty_50 : _GEN_561; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_563 = 8'h33 == req_index ? dirty_51 : _GEN_562; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_564 = 8'h34 == req_index ? dirty_52 : _GEN_563; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_565 = 8'h35 == req_index ? dirty_53 : _GEN_564; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_566 = 8'h36 == req_index ? dirty_54 : _GEN_565; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_567 = 8'h37 == req_index ? dirty_55 : _GEN_566; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_568 = 8'h38 == req_index ? dirty_56 : _GEN_567; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_569 = 8'h39 == req_index ? dirty_57 : _GEN_568; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_570 = 8'h3a == req_index ? dirty_58 : _GEN_569; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_571 = 8'h3b == req_index ? dirty_59 : _GEN_570; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_572 = 8'h3c == req_index ? dirty_60 : _GEN_571; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_573 = 8'h3d == req_index ? dirty_61 : _GEN_572; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_574 = 8'h3e == req_index ? dirty_62 : _GEN_573; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_575 = 8'h3f == req_index ? dirty_63 : _GEN_574; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_576 = 8'h40 == req_index ? dirty_64 : _GEN_575; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_577 = 8'h41 == req_index ? dirty_65 : _GEN_576; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_578 = 8'h42 == req_index ? dirty_66 : _GEN_577; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_579 = 8'h43 == req_index ? dirty_67 : _GEN_578; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_580 = 8'h44 == req_index ? dirty_68 : _GEN_579; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_581 = 8'h45 == req_index ? dirty_69 : _GEN_580; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_582 = 8'h46 == req_index ? dirty_70 : _GEN_581; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_583 = 8'h47 == req_index ? dirty_71 : _GEN_582; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_584 = 8'h48 == req_index ? dirty_72 : _GEN_583; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_585 = 8'h49 == req_index ? dirty_73 : _GEN_584; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_586 = 8'h4a == req_index ? dirty_74 : _GEN_585; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_587 = 8'h4b == req_index ? dirty_75 : _GEN_586; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_588 = 8'h4c == req_index ? dirty_76 : _GEN_587; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_589 = 8'h4d == req_index ? dirty_77 : _GEN_588; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_590 = 8'h4e == req_index ? dirty_78 : _GEN_589; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_591 = 8'h4f == req_index ? dirty_79 : _GEN_590; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_592 = 8'h50 == req_index ? dirty_80 : _GEN_591; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_593 = 8'h51 == req_index ? dirty_81 : _GEN_592; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_594 = 8'h52 == req_index ? dirty_82 : _GEN_593; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_595 = 8'h53 == req_index ? dirty_83 : _GEN_594; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_596 = 8'h54 == req_index ? dirty_84 : _GEN_595; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_597 = 8'h55 == req_index ? dirty_85 : _GEN_596; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_598 = 8'h56 == req_index ? dirty_86 : _GEN_597; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_599 = 8'h57 == req_index ? dirty_87 : _GEN_598; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_600 = 8'h58 == req_index ? dirty_88 : _GEN_599; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_601 = 8'h59 == req_index ? dirty_89 : _GEN_600; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_602 = 8'h5a == req_index ? dirty_90 : _GEN_601; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_603 = 8'h5b == req_index ? dirty_91 : _GEN_602; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_604 = 8'h5c == req_index ? dirty_92 : _GEN_603; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_605 = 8'h5d == req_index ? dirty_93 : _GEN_604; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_606 = 8'h5e == req_index ? dirty_94 : _GEN_605; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_607 = 8'h5f == req_index ? dirty_95 : _GEN_606; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_608 = 8'h60 == req_index ? dirty_96 : _GEN_607; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_609 = 8'h61 == req_index ? dirty_97 : _GEN_608; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_610 = 8'h62 == req_index ? dirty_98 : _GEN_609; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_611 = 8'h63 == req_index ? dirty_99 : _GEN_610; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_612 = 8'h64 == req_index ? dirty_100 : _GEN_611; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_613 = 8'h65 == req_index ? dirty_101 : _GEN_612; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_614 = 8'h66 == req_index ? dirty_102 : _GEN_613; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_615 = 8'h67 == req_index ? dirty_103 : _GEN_614; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_616 = 8'h68 == req_index ? dirty_104 : _GEN_615; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_617 = 8'h69 == req_index ? dirty_105 : _GEN_616; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_618 = 8'h6a == req_index ? dirty_106 : _GEN_617; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_619 = 8'h6b == req_index ? dirty_107 : _GEN_618; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_620 = 8'h6c == req_index ? dirty_108 : _GEN_619; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_621 = 8'h6d == req_index ? dirty_109 : _GEN_620; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_622 = 8'h6e == req_index ? dirty_110 : _GEN_621; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_623 = 8'h6f == req_index ? dirty_111 : _GEN_622; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_624 = 8'h70 == req_index ? dirty_112 : _GEN_623; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_625 = 8'h71 == req_index ? dirty_113 : _GEN_624; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_626 = 8'h72 == req_index ? dirty_114 : _GEN_625; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_627 = 8'h73 == req_index ? dirty_115 : _GEN_626; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_628 = 8'h74 == req_index ? dirty_116 : _GEN_627; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_629 = 8'h75 == req_index ? dirty_117 : _GEN_628; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_630 = 8'h76 == req_index ? dirty_118 : _GEN_629; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_631 = 8'h77 == req_index ? dirty_119 : _GEN_630; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_632 = 8'h78 == req_index ? dirty_120 : _GEN_631; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_633 = 8'h79 == req_index ? dirty_121 : _GEN_632; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_634 = 8'h7a == req_index ? dirty_122 : _GEN_633; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_635 = 8'h7b == req_index ? dirty_123 : _GEN_634; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_636 = 8'h7c == req_index ? dirty_124 : _GEN_635; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_637 = 8'h7d == req_index ? dirty_125 : _GEN_636; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_638 = 8'h7e == req_index ? dirty_126 : _GEN_637; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_639 = 8'h7f == req_index ? dirty_127 : _GEN_638; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_640 = 8'h80 == req_index ? dirty_128 : _GEN_639; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_641 = 8'h81 == req_index ? dirty_129 : _GEN_640; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_642 = 8'h82 == req_index ? dirty_130 : _GEN_641; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_643 = 8'h83 == req_index ? dirty_131 : _GEN_642; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_644 = 8'h84 == req_index ? dirty_132 : _GEN_643; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_645 = 8'h85 == req_index ? dirty_133 : _GEN_644; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_646 = 8'h86 == req_index ? dirty_134 : _GEN_645; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_647 = 8'h87 == req_index ? dirty_135 : _GEN_646; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_648 = 8'h88 == req_index ? dirty_136 : _GEN_647; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_649 = 8'h89 == req_index ? dirty_137 : _GEN_648; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_650 = 8'h8a == req_index ? dirty_138 : _GEN_649; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_651 = 8'h8b == req_index ? dirty_139 : _GEN_650; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_652 = 8'h8c == req_index ? dirty_140 : _GEN_651; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_653 = 8'h8d == req_index ? dirty_141 : _GEN_652; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_654 = 8'h8e == req_index ? dirty_142 : _GEN_653; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_655 = 8'h8f == req_index ? dirty_143 : _GEN_654; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_656 = 8'h90 == req_index ? dirty_144 : _GEN_655; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_657 = 8'h91 == req_index ? dirty_145 : _GEN_656; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_658 = 8'h92 == req_index ? dirty_146 : _GEN_657; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_659 = 8'h93 == req_index ? dirty_147 : _GEN_658; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_660 = 8'h94 == req_index ? dirty_148 : _GEN_659; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_661 = 8'h95 == req_index ? dirty_149 : _GEN_660; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_662 = 8'h96 == req_index ? dirty_150 : _GEN_661; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_663 = 8'h97 == req_index ? dirty_151 : _GEN_662; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_664 = 8'h98 == req_index ? dirty_152 : _GEN_663; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_665 = 8'h99 == req_index ? dirty_153 : _GEN_664; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_666 = 8'h9a == req_index ? dirty_154 : _GEN_665; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_667 = 8'h9b == req_index ? dirty_155 : _GEN_666; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_668 = 8'h9c == req_index ? dirty_156 : _GEN_667; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_669 = 8'h9d == req_index ? dirty_157 : _GEN_668; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_670 = 8'h9e == req_index ? dirty_158 : _GEN_669; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_671 = 8'h9f == req_index ? dirty_159 : _GEN_670; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_672 = 8'ha0 == req_index ? dirty_160 : _GEN_671; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_673 = 8'ha1 == req_index ? dirty_161 : _GEN_672; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_674 = 8'ha2 == req_index ? dirty_162 : _GEN_673; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_675 = 8'ha3 == req_index ? dirty_163 : _GEN_674; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_676 = 8'ha4 == req_index ? dirty_164 : _GEN_675; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_677 = 8'ha5 == req_index ? dirty_165 : _GEN_676; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_678 = 8'ha6 == req_index ? dirty_166 : _GEN_677; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_679 = 8'ha7 == req_index ? dirty_167 : _GEN_678; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_680 = 8'ha8 == req_index ? dirty_168 : _GEN_679; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_681 = 8'ha9 == req_index ? dirty_169 : _GEN_680; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_682 = 8'haa == req_index ? dirty_170 : _GEN_681; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_683 = 8'hab == req_index ? dirty_171 : _GEN_682; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_684 = 8'hac == req_index ? dirty_172 : _GEN_683; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_685 = 8'had == req_index ? dirty_173 : _GEN_684; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_686 = 8'hae == req_index ? dirty_174 : _GEN_685; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_687 = 8'haf == req_index ? dirty_175 : _GEN_686; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_688 = 8'hb0 == req_index ? dirty_176 : _GEN_687; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_689 = 8'hb1 == req_index ? dirty_177 : _GEN_688; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_690 = 8'hb2 == req_index ? dirty_178 : _GEN_689; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_691 = 8'hb3 == req_index ? dirty_179 : _GEN_690; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_692 = 8'hb4 == req_index ? dirty_180 : _GEN_691; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_693 = 8'hb5 == req_index ? dirty_181 : _GEN_692; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_694 = 8'hb6 == req_index ? dirty_182 : _GEN_693; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_695 = 8'hb7 == req_index ? dirty_183 : _GEN_694; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_696 = 8'hb8 == req_index ? dirty_184 : _GEN_695; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_697 = 8'hb9 == req_index ? dirty_185 : _GEN_696; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_698 = 8'hba == req_index ? dirty_186 : _GEN_697; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_699 = 8'hbb == req_index ? dirty_187 : _GEN_698; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_700 = 8'hbc == req_index ? dirty_188 : _GEN_699; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_701 = 8'hbd == req_index ? dirty_189 : _GEN_700; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_702 = 8'hbe == req_index ? dirty_190 : _GEN_701; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_703 = 8'hbf == req_index ? dirty_191 : _GEN_702; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_704 = 8'hc0 == req_index ? dirty_192 : _GEN_703; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_705 = 8'hc1 == req_index ? dirty_193 : _GEN_704; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_706 = 8'hc2 == req_index ? dirty_194 : _GEN_705; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_707 = 8'hc3 == req_index ? dirty_195 : _GEN_706; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_708 = 8'hc4 == req_index ? dirty_196 : _GEN_707; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_709 = 8'hc5 == req_index ? dirty_197 : _GEN_708; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_710 = 8'hc6 == req_index ? dirty_198 : _GEN_709; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_711 = 8'hc7 == req_index ? dirty_199 : _GEN_710; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_712 = 8'hc8 == req_index ? dirty_200 : _GEN_711; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_713 = 8'hc9 == req_index ? dirty_201 : _GEN_712; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_714 = 8'hca == req_index ? dirty_202 : _GEN_713; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_715 = 8'hcb == req_index ? dirty_203 : _GEN_714; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_716 = 8'hcc == req_index ? dirty_204 : _GEN_715; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_717 = 8'hcd == req_index ? dirty_205 : _GEN_716; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_718 = 8'hce == req_index ? dirty_206 : _GEN_717; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_719 = 8'hcf == req_index ? dirty_207 : _GEN_718; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_720 = 8'hd0 == req_index ? dirty_208 : _GEN_719; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_721 = 8'hd1 == req_index ? dirty_209 : _GEN_720; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_722 = 8'hd2 == req_index ? dirty_210 : _GEN_721; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_723 = 8'hd3 == req_index ? dirty_211 : _GEN_722; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_724 = 8'hd4 == req_index ? dirty_212 : _GEN_723; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_725 = 8'hd5 == req_index ? dirty_213 : _GEN_724; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_726 = 8'hd6 == req_index ? dirty_214 : _GEN_725; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_727 = 8'hd7 == req_index ? dirty_215 : _GEN_726; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_728 = 8'hd8 == req_index ? dirty_216 : _GEN_727; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_729 = 8'hd9 == req_index ? dirty_217 : _GEN_728; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_730 = 8'hda == req_index ? dirty_218 : _GEN_729; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_731 = 8'hdb == req_index ? dirty_219 : _GEN_730; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_732 = 8'hdc == req_index ? dirty_220 : _GEN_731; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_733 = 8'hdd == req_index ? dirty_221 : _GEN_732; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_734 = 8'hde == req_index ? dirty_222 : _GEN_733; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_735 = 8'hdf == req_index ? dirty_223 : _GEN_734; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_736 = 8'he0 == req_index ? dirty_224 : _GEN_735; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_737 = 8'he1 == req_index ? dirty_225 : _GEN_736; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_738 = 8'he2 == req_index ? dirty_226 : _GEN_737; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_739 = 8'he3 == req_index ? dirty_227 : _GEN_738; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_740 = 8'he4 == req_index ? dirty_228 : _GEN_739; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_741 = 8'he5 == req_index ? dirty_229 : _GEN_740; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_742 = 8'he6 == req_index ? dirty_230 : _GEN_741; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_743 = 8'he7 == req_index ? dirty_231 : _GEN_742; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_744 = 8'he8 == req_index ? dirty_232 : _GEN_743; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_745 = 8'he9 == req_index ? dirty_233 : _GEN_744; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_746 = 8'hea == req_index ? dirty_234 : _GEN_745; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_747 = 8'heb == req_index ? dirty_235 : _GEN_746; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_748 = 8'hec == req_index ? dirty_236 : _GEN_747; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_749 = 8'hed == req_index ? dirty_237 : _GEN_748; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_750 = 8'hee == req_index ? dirty_238 : _GEN_749; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_751 = 8'hef == req_index ? dirty_239 : _GEN_750; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_752 = 8'hf0 == req_index ? dirty_240 : _GEN_751; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_753 = 8'hf1 == req_index ? dirty_241 : _GEN_752; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_754 = 8'hf2 == req_index ? dirty_242 : _GEN_753; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_755 = 8'hf3 == req_index ? dirty_243 : _GEN_754; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_756 = 8'hf4 == req_index ? dirty_244 : _GEN_755; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_757 = 8'hf5 == req_index ? dirty_245 : _GEN_756; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_758 = 8'hf6 == req_index ? dirty_246 : _GEN_757; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_759 = 8'hf7 == req_index ? dirty_247 : _GEN_758; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_760 = 8'hf8 == req_index ? dirty_248 : _GEN_759; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_761 = 8'hf9 == req_index ? dirty_249 : _GEN_760; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_762 = 8'hfa == req_index ? dirty_250 : _GEN_761; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_763 = 8'hfb == req_index ? dirty_251 : _GEN_762; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_764 = 8'hfc == req_index ? dirty_252 : _GEN_763; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_765 = 8'hfd == req_index ? dirty_253 : _GEN_764; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_766 = 8'hfe == req_index ? dirty_254 : _GEN_765; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  _GEN_767 = 8'hff == req_index ? dirty_255 : _GEN_766; // @[Dcache.scala 35:38 Dcache.scala 35:38]
  wire  cache_dirty = _GEN_767 & _cache_hit_T_2; // @[Dcache.scala 35:38]
  reg  data_ready; // @[Dcache.scala 46:28]
  wire [127:0] cache_data_out = req_Q; // @[Dcache.scala 37:28 Dcache.scala 224:18]
  wire [63:0] valid_rdata = req_offset[3] ? cache_data_out[127:64] : cache_data_out[63:0]; // @[Dcache.scala 48:24]
  wire [7:0] _valid_strb_T_1 = 8'h1 == io_dmem_data_strb ? 8'hff : 8'h0; // @[Mux.scala 80:57]
  wire [15:0] _valid_strb_T_3 = 8'h2 == io_dmem_data_strb ? 16'hff00 : {{8'd0}, _valid_strb_T_1}; // @[Mux.scala 80:57]
  wire [23:0] _valid_strb_T_5 = 8'h4 == io_dmem_data_strb ? 24'hff0000 : {{8'd0}, _valid_strb_T_3}; // @[Mux.scala 80:57]
  wire [31:0] _valid_strb_T_7 = 8'h8 == io_dmem_data_strb ? 32'hff000000 : {{8'd0}, _valid_strb_T_5}; // @[Mux.scala 80:57]
  wire [39:0] _valid_strb_T_9 = 8'h10 == io_dmem_data_strb ? 40'hff00000000 : {{8'd0}, _valid_strb_T_7}; // @[Mux.scala 80:57]
  wire [47:0] _valid_strb_T_11 = 8'h20 == io_dmem_data_strb ? 48'hff0000000000 : {{8'd0}, _valid_strb_T_9}; // @[Mux.scala 80:57]
  wire [55:0] _valid_strb_T_13 = 8'h40 == io_dmem_data_strb ? 56'hff000000000000 : {{8'd0}, _valid_strb_T_11}; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_15 = 8'h80 == io_dmem_data_strb ? 64'hff00000000000000 : {{8'd0}, _valid_strb_T_13}; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_17 = 8'h3 == io_dmem_data_strb ? 64'hffff : _valid_strb_T_15; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_19 = 8'hc == io_dmem_data_strb ? 64'hffff0000 : _valid_strb_T_17; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_21 = 8'h30 == io_dmem_data_strb ? 64'hffff00000000 : _valid_strb_T_19; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_23 = 8'hc0 == io_dmem_data_strb ? 64'hffff000000000000 : _valid_strb_T_21; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_25 = 8'hf == io_dmem_data_strb ? 64'hffffffff : _valid_strb_T_23; // @[Mux.scala 80:57]
  wire [63:0] _valid_strb_T_27 = 8'hf0 == io_dmem_data_strb ? 64'hffffffff00000000 : _valid_strb_T_25; // @[Mux.scala 80:57]
  wire [63:0] valid_strb = 8'hff == io_dmem_data_strb ? 64'hffffffffffffffff : _valid_strb_T_27; // @[Mux.scala 80:57]
  wire [63:0] valid_data = req_offset[3] ? io_out_data_read[127:64] : io_out_data_read[63:0]; // @[Dcache.scala 67:24]
  wire [55:0] valid_wdata_hi = valid_data[63:8]; // @[Dcache.scala 70:47]
  wire [7:0] valid_wdata_lo = io_dmem_data_write[7:0]; // @[Dcache.scala 70:69]
  wire [63:0] _valid_wdata_T_1 = {valid_wdata_hi,valid_wdata_lo}; // @[Cat.scala 30:58]
  wire [47:0] valid_wdata_hi_hi = valid_data[63:16]; // @[Dcache.scala 71:47]
  wire [7:0] valid_wdata_hi_lo = io_dmem_data_write[15:8]; // @[Dcache.scala 71:69]
  wire [7:0] valid_wdata_lo_1 = valid_data[7:0]; // @[Dcache.scala 71:88]
  wire [63:0] _valid_wdata_T_2 = {valid_wdata_hi_hi,valid_wdata_hi_lo,valid_wdata_lo_1}; // @[Cat.scala 30:58]
  wire [39:0] valid_wdata_hi_hi_1 = valid_data[63:24]; // @[Dcache.scala 72:47]
  wire [7:0] valid_wdata_hi_lo_1 = io_dmem_data_write[23:16]; // @[Dcache.scala 72:69]
  wire [15:0] valid_wdata_lo_2 = valid_data[15:0]; // @[Dcache.scala 72:88]
  wire [63:0] _valid_wdata_T_3 = {valid_wdata_hi_hi_1,valid_wdata_hi_lo_1,valid_wdata_lo_2}; // @[Cat.scala 30:58]
  wire [31:0] valid_wdata_hi_hi_2 = valid_data[63:32]; // @[Dcache.scala 73:47]
  wire [7:0] valid_wdata_hi_lo_2 = io_dmem_data_write[31:24]; // @[Dcache.scala 73:69]
  wire [23:0] valid_wdata_lo_3 = valid_data[23:0]; // @[Dcache.scala 73:88]
  wire [63:0] _valid_wdata_T_4 = {valid_wdata_hi_hi_2,valid_wdata_hi_lo_2,valid_wdata_lo_3}; // @[Cat.scala 30:58]
  wire [23:0] valid_wdata_hi_hi_3 = valid_data[63:40]; // @[Dcache.scala 74:47]
  wire [7:0] valid_wdata_hi_lo_3 = io_dmem_data_write[39:32]; // @[Dcache.scala 74:69]
  wire [31:0] valid_wdata_lo_4 = valid_data[31:0]; // @[Dcache.scala 74:88]
  wire [63:0] _valid_wdata_T_5 = {valid_wdata_hi_hi_3,valid_wdata_hi_lo_3,valid_wdata_lo_4}; // @[Cat.scala 30:58]
  wire [15:0] valid_wdata_hi_hi_4 = valid_data[63:48]; // @[Dcache.scala 75:47]
  wire [7:0] valid_wdata_hi_lo_4 = io_dmem_data_write[47:40]; // @[Dcache.scala 75:69]
  wire [39:0] valid_wdata_lo_5 = valid_data[39:0]; // @[Dcache.scala 75:88]
  wire [63:0] _valid_wdata_T_6 = {valid_wdata_hi_hi_4,valid_wdata_hi_lo_4,valid_wdata_lo_5}; // @[Cat.scala 30:58]
  wire [7:0] valid_wdata_hi_hi_5 = valid_data[63:56]; // @[Dcache.scala 76:47]
  wire [7:0] valid_wdata_hi_lo_5 = io_dmem_data_write[55:48]; // @[Dcache.scala 76:69]
  wire [47:0] valid_wdata_lo_6 = valid_data[47:0]; // @[Dcache.scala 76:88]
  wire [63:0] _valid_wdata_T_7 = {valid_wdata_hi_hi_5,valid_wdata_hi_lo_5,valid_wdata_lo_6}; // @[Cat.scala 30:58]
  wire [7:0] valid_wdata_hi_7 = io_dmem_data_write[63:56]; // @[Dcache.scala 77:50]
  wire [55:0] valid_wdata_lo_7 = valid_data[55:0]; // @[Dcache.scala 77:69]
  wire [63:0] _valid_wdata_T_8 = {valid_wdata_hi_7,valid_wdata_lo_7}; // @[Cat.scala 30:58]
  wire [63:0] _valid_wdata_T_10 = 3'h1 == req_offset[2:0] ? _valid_wdata_T_2 : _valid_wdata_T_1; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_12 = 3'h2 == req_offset[2:0] ? _valid_wdata_T_3 : _valid_wdata_T_10; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_14 = 3'h3 == req_offset[2:0] ? _valid_wdata_T_4 : _valid_wdata_T_12; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_16 = 3'h4 == req_offset[2:0] ? _valid_wdata_T_5 : _valid_wdata_T_14; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_18 = 3'h5 == req_offset[2:0] ? _valid_wdata_T_6 : _valid_wdata_T_16; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_20 = 3'h6 == req_offset[2:0] ? _valid_wdata_T_7 : _valid_wdata_T_18; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_22 = 3'h7 == req_offset[2:0] ? _valid_wdata_T_8 : _valid_wdata_T_20; // @[Mux.scala 80:57]
  wire [15:0] valid_wdata_lo_8 = io_dmem_data_write[15:0]; // @[Dcache.scala 80:68]
  wire [63:0] _valid_wdata_T_24 = {valid_wdata_hi_hi,valid_wdata_lo_8}; // @[Cat.scala 30:58]
  wire [15:0] valid_wdata_hi_lo_6 = io_dmem_data_write[31:16]; // @[Dcache.scala 81:68]
  wire [63:0] _valid_wdata_T_25 = {valid_wdata_hi_hi_2,valid_wdata_hi_lo_6,valid_wdata_lo_2}; // @[Cat.scala 30:58]
  wire [15:0] valid_wdata_hi_lo_7 = io_dmem_data_write[47:32]; // @[Dcache.scala 82:68]
  wire [63:0] _valid_wdata_T_26 = {valid_wdata_hi_hi_4,valid_wdata_hi_lo_7,valid_wdata_lo_4}; // @[Cat.scala 30:58]
  wire [15:0] valid_wdata_hi_11 = io_dmem_data_write[63:48]; // @[Dcache.scala 83:49]
  wire [63:0] _valid_wdata_T_27 = {valid_wdata_hi_11,valid_wdata_lo_6}; // @[Cat.scala 30:58]
  wire [63:0] _valid_wdata_T_29 = 2'h1 == req_offset[2:1] ? _valid_wdata_T_25 : _valid_wdata_T_24; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_31 = 2'h2 == req_offset[2:1] ? _valid_wdata_T_26 : _valid_wdata_T_29; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_33 = 2'h3 == req_offset[2:1] ? _valid_wdata_T_27 : _valid_wdata_T_31; // @[Mux.scala 80:57]
  wire [31:0] valid_wdata_lo_12 = io_dmem_data_write[31:0]; // @[Dcache.scala 86:67]
  wire [63:0] _valid_wdata_T_35 = {valid_wdata_hi_hi_2,valid_wdata_lo_12}; // @[Cat.scala 30:58]
  wire [31:0] valid_wdata_hi_13 = io_dmem_data_write[63:32]; // @[Dcache.scala 87:48]
  wire [63:0] _valid_wdata_T_36 = {valid_wdata_hi_13,valid_wdata_lo_4}; // @[Cat.scala 30:58]
  wire [63:0] _valid_wdata_T_38 = req_offset[2] ? _valid_wdata_T_36 : _valid_wdata_T_35; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_40 = 2'h1 == io_dmem_data_size ? _valid_wdata_T_33 : _valid_wdata_T_22; // @[Mux.scala 80:57]
  wire [63:0] _valid_wdata_T_42 = 2'h2 == io_dmem_data_size ? _valid_wdata_T_38 : _valid_wdata_T_40; // @[Mux.scala 80:57]
  wire [63:0] valid_wdata = 2'h3 == io_dmem_data_size ? io_dmem_data_write : _valid_wdata_T_42; // @[Mux.scala 80:57]
  wire [7:0] data_read_lo = valid_rdata[7:0]; // @[Dcache.scala 94:53]
  wire [8:0] _data_read_T_1 = {1'h0,data_read_lo}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_1 = valid_rdata[15:8]; // @[Dcache.scala 95:53]
  wire [8:0] _data_read_T_2 = {1'h0,data_read_lo_1}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_2 = valid_rdata[23:16]; // @[Dcache.scala 96:53]
  wire [8:0] _data_read_T_3 = {1'h0,data_read_lo_2}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_3 = valid_rdata[31:24]; // @[Dcache.scala 97:53]
  wire [8:0] _data_read_T_4 = {1'h0,data_read_lo_3}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_4 = valid_rdata[39:32]; // @[Dcache.scala 98:53]
  wire [8:0] _data_read_T_5 = {1'h0,data_read_lo_4}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_5 = valid_rdata[47:40]; // @[Dcache.scala 99:53]
  wire [8:0] _data_read_T_6 = {1'h0,data_read_lo_5}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_6 = valid_rdata[55:48]; // @[Dcache.scala 100:53]
  wire [8:0] _data_read_T_7 = {1'h0,data_read_lo_6}; // @[Cat.scala 30:58]
  wire [7:0] data_read_lo_7 = valid_rdata[63:56]; // @[Dcache.scala 101:53]
  wire [8:0] _data_read_T_8 = {1'h0,data_read_lo_7}; // @[Cat.scala 30:58]
  wire [8:0] _data_read_T_10 = 3'h1 == req_offset[2:0] ? _data_read_T_2 : _data_read_T_1; // @[Mux.scala 80:57]
  wire [8:0] _data_read_T_12 = 3'h2 == req_offset[2:0] ? _data_read_T_3 : _data_read_T_10; // @[Mux.scala 80:57]
  wire [8:0] _data_read_T_14 = 3'h3 == req_offset[2:0] ? _data_read_T_4 : _data_read_T_12; // @[Mux.scala 80:57]
  wire [8:0] _data_read_T_16 = 3'h4 == req_offset[2:0] ? _data_read_T_5 : _data_read_T_14; // @[Mux.scala 80:57]
  wire [8:0] _data_read_T_18 = 3'h5 == req_offset[2:0] ? _data_read_T_6 : _data_read_T_16; // @[Mux.scala 80:57]
  wire [8:0] _data_read_T_20 = 3'h6 == req_offset[2:0] ? _data_read_T_7 : _data_read_T_18; // @[Mux.scala 80:57]
  wire [8:0] _data_read_T_22 = 3'h7 == req_offset[2:0] ? _data_read_T_8 : _data_read_T_20; // @[Mux.scala 80:57]
  wire [15:0] data_read_lo_8 = valid_rdata[15:0]; // @[Dcache.scala 104:52]
  wire [16:0] _data_read_T_24 = {1'h0,data_read_lo_8}; // @[Cat.scala 30:58]
  wire [15:0] data_read_lo_9 = valid_rdata[31:16]; // @[Dcache.scala 105:52]
  wire [16:0] _data_read_T_25 = {1'h0,data_read_lo_9}; // @[Cat.scala 30:58]
  wire [15:0] data_read_lo_10 = valid_rdata[47:32]; // @[Dcache.scala 106:52]
  wire [16:0] _data_read_T_26 = {1'h0,data_read_lo_10}; // @[Cat.scala 30:58]
  wire [15:0] data_read_lo_11 = valid_rdata[63:48]; // @[Dcache.scala 107:52]
  wire [16:0] _data_read_T_27 = {1'h0,data_read_lo_11}; // @[Cat.scala 30:58]
  wire [16:0] _data_read_T_29 = 2'h1 == req_offset[2:1] ? _data_read_T_25 : _data_read_T_24; // @[Mux.scala 80:57]
  wire [16:0] _data_read_T_31 = 2'h2 == req_offset[2:1] ? _data_read_T_26 : _data_read_T_29; // @[Mux.scala 80:57]
  wire [16:0] _data_read_T_33 = 2'h3 == req_offset[2:1] ? _data_read_T_27 : _data_read_T_31; // @[Mux.scala 80:57]
  wire [31:0] data_read_lo_12 = valid_rdata[31:0]; // @[Dcache.scala 110:51]
  wire [32:0] _data_read_T_35 = {1'h0,data_read_lo_12}; // @[Cat.scala 30:58]
  wire [31:0] data_read_lo_13 = valid_rdata[63:32]; // @[Dcache.scala 111:51]
  wire [32:0] _data_read_T_36 = {1'h0,data_read_lo_13}; // @[Cat.scala 30:58]
  wire [32:0] _data_read_T_38 = req_offset[2] ? _data_read_T_36 : _data_read_T_35; // @[Mux.scala 80:57]
  wire [16:0] _data_read_T_40 = 2'h1 == io_dmem_data_size ? _data_read_T_33 : {{8'd0}, _data_read_T_22}; // @[Mux.scala 80:57]
  wire [32:0] _data_read_T_42 = 2'h2 == io_dmem_data_size ? _data_read_T_38 : {{16'd0}, _data_read_T_40}; // @[Mux.scala 80:57]
  reg  cache_fill; // @[Dcache.scala 116:28]
  reg  cache_wen; // @[Dcache.scala 117:28]
  reg [127:0] cache_wdata; // @[Dcache.scala 118:28]
  reg [127:0] cache_strb; // @[Dcache.scala 119:28]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _GEN_769 = 8'h0 == req_index | valid_0; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_770 = 8'h1 == req_index | valid_1; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_771 = 8'h2 == req_index | valid_2; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_772 = 8'h3 == req_index | valid_3; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_773 = 8'h4 == req_index | valid_4; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_774 = 8'h5 == req_index | valid_5; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_775 = 8'h6 == req_index | valid_6; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_776 = 8'h7 == req_index | valid_7; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_777 = 8'h8 == req_index | valid_8; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_778 = 8'h9 == req_index | valid_9; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_779 = 8'ha == req_index | valid_10; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_780 = 8'hb == req_index | valid_11; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_781 = 8'hc == req_index | valid_12; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_782 = 8'hd == req_index | valid_13; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_783 = 8'he == req_index | valid_14; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_784 = 8'hf == req_index | valid_15; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_785 = 8'h10 == req_index | valid_16; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_786 = 8'h11 == req_index | valid_17; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_787 = 8'h12 == req_index | valid_18; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_788 = 8'h13 == req_index | valid_19; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_789 = 8'h14 == req_index | valid_20; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_790 = 8'h15 == req_index | valid_21; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_791 = 8'h16 == req_index | valid_22; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_792 = 8'h17 == req_index | valid_23; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_793 = 8'h18 == req_index | valid_24; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_794 = 8'h19 == req_index | valid_25; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_795 = 8'h1a == req_index | valid_26; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_796 = 8'h1b == req_index | valid_27; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_797 = 8'h1c == req_index | valid_28; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_798 = 8'h1d == req_index | valid_29; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_799 = 8'h1e == req_index | valid_30; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_800 = 8'h1f == req_index | valid_31; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_801 = 8'h20 == req_index | valid_32; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_802 = 8'h21 == req_index | valid_33; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_803 = 8'h22 == req_index | valid_34; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_804 = 8'h23 == req_index | valid_35; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_805 = 8'h24 == req_index | valid_36; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_806 = 8'h25 == req_index | valid_37; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_807 = 8'h26 == req_index | valid_38; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_808 = 8'h27 == req_index | valid_39; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_809 = 8'h28 == req_index | valid_40; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_810 = 8'h29 == req_index | valid_41; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_811 = 8'h2a == req_index | valid_42; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_812 = 8'h2b == req_index | valid_43; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_813 = 8'h2c == req_index | valid_44; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_814 = 8'h2d == req_index | valid_45; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_815 = 8'h2e == req_index | valid_46; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_816 = 8'h2f == req_index | valid_47; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_817 = 8'h30 == req_index | valid_48; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_818 = 8'h31 == req_index | valid_49; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_819 = 8'h32 == req_index | valid_50; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_820 = 8'h33 == req_index | valid_51; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_821 = 8'h34 == req_index | valid_52; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_822 = 8'h35 == req_index | valid_53; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_823 = 8'h36 == req_index | valid_54; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_824 = 8'h37 == req_index | valid_55; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_825 = 8'h38 == req_index | valid_56; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_826 = 8'h39 == req_index | valid_57; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_827 = 8'h3a == req_index | valid_58; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_828 = 8'h3b == req_index | valid_59; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_829 = 8'h3c == req_index | valid_60; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_830 = 8'h3d == req_index | valid_61; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_831 = 8'h3e == req_index | valid_62; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_832 = 8'h3f == req_index | valid_63; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_833 = 8'h40 == req_index | valid_64; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_834 = 8'h41 == req_index | valid_65; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_835 = 8'h42 == req_index | valid_66; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_836 = 8'h43 == req_index | valid_67; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_837 = 8'h44 == req_index | valid_68; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_838 = 8'h45 == req_index | valid_69; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_839 = 8'h46 == req_index | valid_70; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_840 = 8'h47 == req_index | valid_71; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_841 = 8'h48 == req_index | valid_72; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_842 = 8'h49 == req_index | valid_73; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_843 = 8'h4a == req_index | valid_74; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_844 = 8'h4b == req_index | valid_75; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_845 = 8'h4c == req_index | valid_76; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_846 = 8'h4d == req_index | valid_77; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_847 = 8'h4e == req_index | valid_78; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_848 = 8'h4f == req_index | valid_79; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_849 = 8'h50 == req_index | valid_80; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_850 = 8'h51 == req_index | valid_81; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_851 = 8'h52 == req_index | valid_82; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_852 = 8'h53 == req_index | valid_83; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_853 = 8'h54 == req_index | valid_84; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_854 = 8'h55 == req_index | valid_85; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_855 = 8'h56 == req_index | valid_86; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_856 = 8'h57 == req_index | valid_87; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_857 = 8'h58 == req_index | valid_88; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_858 = 8'h59 == req_index | valid_89; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_859 = 8'h5a == req_index | valid_90; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_860 = 8'h5b == req_index | valid_91; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_861 = 8'h5c == req_index | valid_92; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_862 = 8'h5d == req_index | valid_93; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_863 = 8'h5e == req_index | valid_94; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_864 = 8'h5f == req_index | valid_95; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_865 = 8'h60 == req_index | valid_96; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_866 = 8'h61 == req_index | valid_97; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_867 = 8'h62 == req_index | valid_98; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_868 = 8'h63 == req_index | valid_99; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_869 = 8'h64 == req_index | valid_100; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_870 = 8'h65 == req_index | valid_101; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_871 = 8'h66 == req_index | valid_102; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_872 = 8'h67 == req_index | valid_103; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_873 = 8'h68 == req_index | valid_104; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_874 = 8'h69 == req_index | valid_105; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_875 = 8'h6a == req_index | valid_106; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_876 = 8'h6b == req_index | valid_107; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_877 = 8'h6c == req_index | valid_108; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_878 = 8'h6d == req_index | valid_109; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_879 = 8'h6e == req_index | valid_110; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_880 = 8'h6f == req_index | valid_111; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_881 = 8'h70 == req_index | valid_112; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_882 = 8'h71 == req_index | valid_113; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_883 = 8'h72 == req_index | valid_114; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_884 = 8'h73 == req_index | valid_115; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_885 = 8'h74 == req_index | valid_116; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_886 = 8'h75 == req_index | valid_117; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_887 = 8'h76 == req_index | valid_118; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_888 = 8'h77 == req_index | valid_119; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_889 = 8'h78 == req_index | valid_120; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_890 = 8'h79 == req_index | valid_121; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_891 = 8'h7a == req_index | valid_122; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_892 = 8'h7b == req_index | valid_123; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_893 = 8'h7c == req_index | valid_124; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_894 = 8'h7d == req_index | valid_125; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_895 = 8'h7e == req_index | valid_126; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_896 = 8'h7f == req_index | valid_127; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_897 = 8'h80 == req_index | valid_128; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_898 = 8'h81 == req_index | valid_129; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_899 = 8'h82 == req_index | valid_130; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_900 = 8'h83 == req_index | valid_131; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_901 = 8'h84 == req_index | valid_132; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_902 = 8'h85 == req_index | valid_133; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_903 = 8'h86 == req_index | valid_134; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_904 = 8'h87 == req_index | valid_135; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_905 = 8'h88 == req_index | valid_136; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_906 = 8'h89 == req_index | valid_137; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_907 = 8'h8a == req_index | valid_138; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_908 = 8'h8b == req_index | valid_139; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_909 = 8'h8c == req_index | valid_140; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_910 = 8'h8d == req_index | valid_141; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_911 = 8'h8e == req_index | valid_142; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_912 = 8'h8f == req_index | valid_143; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_913 = 8'h90 == req_index | valid_144; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_914 = 8'h91 == req_index | valid_145; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_915 = 8'h92 == req_index | valid_146; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_916 = 8'h93 == req_index | valid_147; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_917 = 8'h94 == req_index | valid_148; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_918 = 8'h95 == req_index | valid_149; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_919 = 8'h96 == req_index | valid_150; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_920 = 8'h97 == req_index | valid_151; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_921 = 8'h98 == req_index | valid_152; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_922 = 8'h99 == req_index | valid_153; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_923 = 8'h9a == req_index | valid_154; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_924 = 8'h9b == req_index | valid_155; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_925 = 8'h9c == req_index | valid_156; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_926 = 8'h9d == req_index | valid_157; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_927 = 8'h9e == req_index | valid_158; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_928 = 8'h9f == req_index | valid_159; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_929 = 8'ha0 == req_index | valid_160; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_930 = 8'ha1 == req_index | valid_161; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_931 = 8'ha2 == req_index | valid_162; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_932 = 8'ha3 == req_index | valid_163; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_933 = 8'ha4 == req_index | valid_164; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_934 = 8'ha5 == req_index | valid_165; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_935 = 8'ha6 == req_index | valid_166; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_936 = 8'ha7 == req_index | valid_167; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_937 = 8'ha8 == req_index | valid_168; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_938 = 8'ha9 == req_index | valid_169; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_939 = 8'haa == req_index | valid_170; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_940 = 8'hab == req_index | valid_171; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_941 = 8'hac == req_index | valid_172; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_942 = 8'had == req_index | valid_173; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_943 = 8'hae == req_index | valid_174; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_944 = 8'haf == req_index | valid_175; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_945 = 8'hb0 == req_index | valid_176; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_946 = 8'hb1 == req_index | valid_177; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_947 = 8'hb2 == req_index | valid_178; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_948 = 8'hb3 == req_index | valid_179; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_949 = 8'hb4 == req_index | valid_180; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_950 = 8'hb5 == req_index | valid_181; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_951 = 8'hb6 == req_index | valid_182; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_952 = 8'hb7 == req_index | valid_183; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_953 = 8'hb8 == req_index | valid_184; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_954 = 8'hb9 == req_index | valid_185; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_955 = 8'hba == req_index | valid_186; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_956 = 8'hbb == req_index | valid_187; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_957 = 8'hbc == req_index | valid_188; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_958 = 8'hbd == req_index | valid_189; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_959 = 8'hbe == req_index | valid_190; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_960 = 8'hbf == req_index | valid_191; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_961 = 8'hc0 == req_index | valid_192; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_962 = 8'hc1 == req_index | valid_193; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_963 = 8'hc2 == req_index | valid_194; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_964 = 8'hc3 == req_index | valid_195; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_965 = 8'hc4 == req_index | valid_196; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_966 = 8'hc5 == req_index | valid_197; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_967 = 8'hc6 == req_index | valid_198; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_968 = 8'hc7 == req_index | valid_199; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_969 = 8'hc8 == req_index | valid_200; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_970 = 8'hc9 == req_index | valid_201; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_971 = 8'hca == req_index | valid_202; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_972 = 8'hcb == req_index | valid_203; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_973 = 8'hcc == req_index | valid_204; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_974 = 8'hcd == req_index | valid_205; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_975 = 8'hce == req_index | valid_206; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_976 = 8'hcf == req_index | valid_207; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_977 = 8'hd0 == req_index | valid_208; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_978 = 8'hd1 == req_index | valid_209; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_979 = 8'hd2 == req_index | valid_210; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_980 = 8'hd3 == req_index | valid_211; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_981 = 8'hd4 == req_index | valid_212; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_982 = 8'hd5 == req_index | valid_213; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_983 = 8'hd6 == req_index | valid_214; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_984 = 8'hd7 == req_index | valid_215; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_985 = 8'hd8 == req_index | valid_216; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_986 = 8'hd9 == req_index | valid_217; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_987 = 8'hda == req_index | valid_218; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_988 = 8'hdb == req_index | valid_219; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_989 = 8'hdc == req_index | valid_220; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_990 = 8'hdd == req_index | valid_221; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_991 = 8'hde == req_index | valid_222; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_992 = 8'hdf == req_index | valid_223; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_993 = 8'he0 == req_index | valid_224; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_994 = 8'he1 == req_index | valid_225; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_995 = 8'he2 == req_index | valid_226; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_996 = 8'he3 == req_index | valid_227; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_997 = 8'he4 == req_index | valid_228; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_998 = 8'he5 == req_index | valid_229; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_999 = 8'he6 == req_index | valid_230; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1000 = 8'he7 == req_index | valid_231; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1001 = 8'he8 == req_index | valid_232; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1002 = 8'he9 == req_index | valid_233; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1003 = 8'hea == req_index | valid_234; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1004 = 8'heb == req_index | valid_235; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1005 = 8'hec == req_index | valid_236; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1006 = 8'hed == req_index | valid_237; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1007 = 8'hee == req_index | valid_238; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1008 = 8'hef == req_index | valid_239; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1009 = 8'hf0 == req_index | valid_240; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1010 = 8'hf1 == req_index | valid_241; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1011 = 8'hf2 == req_index | valid_242; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1012 = 8'hf3 == req_index | valid_243; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1013 = 8'hf4 == req_index | valid_244; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1014 = 8'hf5 == req_index | valid_245; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1015 = 8'hf6 == req_index | valid_246; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1016 = 8'hf7 == req_index | valid_247; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1017 = 8'hf8 == req_index | valid_248; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1018 = 8'hf9 == req_index | valid_249; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1019 = 8'hfa == req_index | valid_250; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1020 = 8'hfb == req_index | valid_251; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1021 = 8'hfc == req_index | valid_252; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1022 = 8'hfd == req_index | valid_253; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1023 = 8'hfe == req_index | valid_254; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire  _GEN_1024 = 8'hff == req_index | valid_255; // @[Dcache.scala 132:27 Dcache.scala 132:27 Dcache.scala 17:24]
  wire [19:0] _GEN_1025 = 8'h0 == req_index ? req_tag : tag_0; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1026 = 8'h1 == req_index ? req_tag : tag_1; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1027 = 8'h2 == req_index ? req_tag : tag_2; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1028 = 8'h3 == req_index ? req_tag : tag_3; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1029 = 8'h4 == req_index ? req_tag : tag_4; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1030 = 8'h5 == req_index ? req_tag : tag_5; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1031 = 8'h6 == req_index ? req_tag : tag_6; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1032 = 8'h7 == req_index ? req_tag : tag_7; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1033 = 8'h8 == req_index ? req_tag : tag_8; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1034 = 8'h9 == req_index ? req_tag : tag_9; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1035 = 8'ha == req_index ? req_tag : tag_10; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1036 = 8'hb == req_index ? req_tag : tag_11; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1037 = 8'hc == req_index ? req_tag : tag_12; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1038 = 8'hd == req_index ? req_tag : tag_13; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1039 = 8'he == req_index ? req_tag : tag_14; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1040 = 8'hf == req_index ? req_tag : tag_15; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1041 = 8'h10 == req_index ? req_tag : tag_16; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1042 = 8'h11 == req_index ? req_tag : tag_17; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1043 = 8'h12 == req_index ? req_tag : tag_18; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1044 = 8'h13 == req_index ? req_tag : tag_19; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1045 = 8'h14 == req_index ? req_tag : tag_20; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1046 = 8'h15 == req_index ? req_tag : tag_21; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1047 = 8'h16 == req_index ? req_tag : tag_22; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1048 = 8'h17 == req_index ? req_tag : tag_23; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1049 = 8'h18 == req_index ? req_tag : tag_24; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1050 = 8'h19 == req_index ? req_tag : tag_25; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1051 = 8'h1a == req_index ? req_tag : tag_26; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1052 = 8'h1b == req_index ? req_tag : tag_27; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1053 = 8'h1c == req_index ? req_tag : tag_28; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1054 = 8'h1d == req_index ? req_tag : tag_29; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1055 = 8'h1e == req_index ? req_tag : tag_30; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1056 = 8'h1f == req_index ? req_tag : tag_31; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1057 = 8'h20 == req_index ? req_tag : tag_32; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1058 = 8'h21 == req_index ? req_tag : tag_33; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1059 = 8'h22 == req_index ? req_tag : tag_34; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1060 = 8'h23 == req_index ? req_tag : tag_35; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1061 = 8'h24 == req_index ? req_tag : tag_36; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1062 = 8'h25 == req_index ? req_tag : tag_37; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1063 = 8'h26 == req_index ? req_tag : tag_38; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1064 = 8'h27 == req_index ? req_tag : tag_39; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1065 = 8'h28 == req_index ? req_tag : tag_40; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1066 = 8'h29 == req_index ? req_tag : tag_41; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1067 = 8'h2a == req_index ? req_tag : tag_42; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1068 = 8'h2b == req_index ? req_tag : tag_43; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1069 = 8'h2c == req_index ? req_tag : tag_44; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1070 = 8'h2d == req_index ? req_tag : tag_45; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1071 = 8'h2e == req_index ? req_tag : tag_46; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1072 = 8'h2f == req_index ? req_tag : tag_47; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1073 = 8'h30 == req_index ? req_tag : tag_48; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1074 = 8'h31 == req_index ? req_tag : tag_49; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1075 = 8'h32 == req_index ? req_tag : tag_50; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1076 = 8'h33 == req_index ? req_tag : tag_51; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1077 = 8'h34 == req_index ? req_tag : tag_52; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1078 = 8'h35 == req_index ? req_tag : tag_53; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1079 = 8'h36 == req_index ? req_tag : tag_54; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1080 = 8'h37 == req_index ? req_tag : tag_55; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1081 = 8'h38 == req_index ? req_tag : tag_56; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1082 = 8'h39 == req_index ? req_tag : tag_57; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1083 = 8'h3a == req_index ? req_tag : tag_58; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1084 = 8'h3b == req_index ? req_tag : tag_59; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1085 = 8'h3c == req_index ? req_tag : tag_60; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1086 = 8'h3d == req_index ? req_tag : tag_61; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1087 = 8'h3e == req_index ? req_tag : tag_62; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1088 = 8'h3f == req_index ? req_tag : tag_63; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1089 = 8'h40 == req_index ? req_tag : tag_64; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1090 = 8'h41 == req_index ? req_tag : tag_65; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1091 = 8'h42 == req_index ? req_tag : tag_66; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1092 = 8'h43 == req_index ? req_tag : tag_67; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1093 = 8'h44 == req_index ? req_tag : tag_68; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1094 = 8'h45 == req_index ? req_tag : tag_69; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1095 = 8'h46 == req_index ? req_tag : tag_70; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1096 = 8'h47 == req_index ? req_tag : tag_71; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1097 = 8'h48 == req_index ? req_tag : tag_72; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1098 = 8'h49 == req_index ? req_tag : tag_73; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1099 = 8'h4a == req_index ? req_tag : tag_74; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1100 = 8'h4b == req_index ? req_tag : tag_75; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1101 = 8'h4c == req_index ? req_tag : tag_76; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1102 = 8'h4d == req_index ? req_tag : tag_77; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1103 = 8'h4e == req_index ? req_tag : tag_78; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1104 = 8'h4f == req_index ? req_tag : tag_79; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1105 = 8'h50 == req_index ? req_tag : tag_80; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1106 = 8'h51 == req_index ? req_tag : tag_81; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1107 = 8'h52 == req_index ? req_tag : tag_82; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1108 = 8'h53 == req_index ? req_tag : tag_83; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1109 = 8'h54 == req_index ? req_tag : tag_84; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1110 = 8'h55 == req_index ? req_tag : tag_85; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1111 = 8'h56 == req_index ? req_tag : tag_86; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1112 = 8'h57 == req_index ? req_tag : tag_87; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1113 = 8'h58 == req_index ? req_tag : tag_88; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1114 = 8'h59 == req_index ? req_tag : tag_89; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1115 = 8'h5a == req_index ? req_tag : tag_90; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1116 = 8'h5b == req_index ? req_tag : tag_91; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1117 = 8'h5c == req_index ? req_tag : tag_92; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1118 = 8'h5d == req_index ? req_tag : tag_93; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1119 = 8'h5e == req_index ? req_tag : tag_94; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1120 = 8'h5f == req_index ? req_tag : tag_95; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1121 = 8'h60 == req_index ? req_tag : tag_96; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1122 = 8'h61 == req_index ? req_tag : tag_97; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1123 = 8'h62 == req_index ? req_tag : tag_98; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1124 = 8'h63 == req_index ? req_tag : tag_99; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1125 = 8'h64 == req_index ? req_tag : tag_100; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1126 = 8'h65 == req_index ? req_tag : tag_101; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1127 = 8'h66 == req_index ? req_tag : tag_102; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1128 = 8'h67 == req_index ? req_tag : tag_103; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1129 = 8'h68 == req_index ? req_tag : tag_104; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1130 = 8'h69 == req_index ? req_tag : tag_105; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1131 = 8'h6a == req_index ? req_tag : tag_106; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1132 = 8'h6b == req_index ? req_tag : tag_107; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1133 = 8'h6c == req_index ? req_tag : tag_108; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1134 = 8'h6d == req_index ? req_tag : tag_109; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1135 = 8'h6e == req_index ? req_tag : tag_110; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1136 = 8'h6f == req_index ? req_tag : tag_111; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1137 = 8'h70 == req_index ? req_tag : tag_112; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1138 = 8'h71 == req_index ? req_tag : tag_113; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1139 = 8'h72 == req_index ? req_tag : tag_114; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1140 = 8'h73 == req_index ? req_tag : tag_115; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1141 = 8'h74 == req_index ? req_tag : tag_116; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1142 = 8'h75 == req_index ? req_tag : tag_117; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1143 = 8'h76 == req_index ? req_tag : tag_118; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1144 = 8'h77 == req_index ? req_tag : tag_119; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1145 = 8'h78 == req_index ? req_tag : tag_120; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1146 = 8'h79 == req_index ? req_tag : tag_121; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1147 = 8'h7a == req_index ? req_tag : tag_122; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1148 = 8'h7b == req_index ? req_tag : tag_123; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1149 = 8'h7c == req_index ? req_tag : tag_124; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1150 = 8'h7d == req_index ? req_tag : tag_125; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1151 = 8'h7e == req_index ? req_tag : tag_126; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1152 = 8'h7f == req_index ? req_tag : tag_127; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1153 = 8'h80 == req_index ? req_tag : tag_128; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1154 = 8'h81 == req_index ? req_tag : tag_129; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1155 = 8'h82 == req_index ? req_tag : tag_130; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1156 = 8'h83 == req_index ? req_tag : tag_131; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1157 = 8'h84 == req_index ? req_tag : tag_132; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1158 = 8'h85 == req_index ? req_tag : tag_133; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1159 = 8'h86 == req_index ? req_tag : tag_134; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1160 = 8'h87 == req_index ? req_tag : tag_135; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1161 = 8'h88 == req_index ? req_tag : tag_136; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1162 = 8'h89 == req_index ? req_tag : tag_137; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1163 = 8'h8a == req_index ? req_tag : tag_138; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1164 = 8'h8b == req_index ? req_tag : tag_139; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1165 = 8'h8c == req_index ? req_tag : tag_140; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1166 = 8'h8d == req_index ? req_tag : tag_141; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1167 = 8'h8e == req_index ? req_tag : tag_142; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1168 = 8'h8f == req_index ? req_tag : tag_143; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1169 = 8'h90 == req_index ? req_tag : tag_144; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1170 = 8'h91 == req_index ? req_tag : tag_145; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1171 = 8'h92 == req_index ? req_tag : tag_146; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1172 = 8'h93 == req_index ? req_tag : tag_147; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1173 = 8'h94 == req_index ? req_tag : tag_148; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1174 = 8'h95 == req_index ? req_tag : tag_149; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1175 = 8'h96 == req_index ? req_tag : tag_150; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1176 = 8'h97 == req_index ? req_tag : tag_151; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1177 = 8'h98 == req_index ? req_tag : tag_152; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1178 = 8'h99 == req_index ? req_tag : tag_153; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1179 = 8'h9a == req_index ? req_tag : tag_154; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1180 = 8'h9b == req_index ? req_tag : tag_155; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1181 = 8'h9c == req_index ? req_tag : tag_156; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1182 = 8'h9d == req_index ? req_tag : tag_157; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1183 = 8'h9e == req_index ? req_tag : tag_158; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1184 = 8'h9f == req_index ? req_tag : tag_159; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1185 = 8'ha0 == req_index ? req_tag : tag_160; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1186 = 8'ha1 == req_index ? req_tag : tag_161; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1187 = 8'ha2 == req_index ? req_tag : tag_162; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1188 = 8'ha3 == req_index ? req_tag : tag_163; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1189 = 8'ha4 == req_index ? req_tag : tag_164; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1190 = 8'ha5 == req_index ? req_tag : tag_165; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1191 = 8'ha6 == req_index ? req_tag : tag_166; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1192 = 8'ha7 == req_index ? req_tag : tag_167; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1193 = 8'ha8 == req_index ? req_tag : tag_168; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1194 = 8'ha9 == req_index ? req_tag : tag_169; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1195 = 8'haa == req_index ? req_tag : tag_170; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1196 = 8'hab == req_index ? req_tag : tag_171; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1197 = 8'hac == req_index ? req_tag : tag_172; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1198 = 8'had == req_index ? req_tag : tag_173; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1199 = 8'hae == req_index ? req_tag : tag_174; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1200 = 8'haf == req_index ? req_tag : tag_175; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1201 = 8'hb0 == req_index ? req_tag : tag_176; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1202 = 8'hb1 == req_index ? req_tag : tag_177; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1203 = 8'hb2 == req_index ? req_tag : tag_178; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1204 = 8'hb3 == req_index ? req_tag : tag_179; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1205 = 8'hb4 == req_index ? req_tag : tag_180; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1206 = 8'hb5 == req_index ? req_tag : tag_181; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1207 = 8'hb6 == req_index ? req_tag : tag_182; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1208 = 8'hb7 == req_index ? req_tag : tag_183; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1209 = 8'hb8 == req_index ? req_tag : tag_184; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1210 = 8'hb9 == req_index ? req_tag : tag_185; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1211 = 8'hba == req_index ? req_tag : tag_186; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1212 = 8'hbb == req_index ? req_tag : tag_187; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1213 = 8'hbc == req_index ? req_tag : tag_188; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1214 = 8'hbd == req_index ? req_tag : tag_189; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1215 = 8'hbe == req_index ? req_tag : tag_190; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1216 = 8'hbf == req_index ? req_tag : tag_191; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1217 = 8'hc0 == req_index ? req_tag : tag_192; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1218 = 8'hc1 == req_index ? req_tag : tag_193; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1219 = 8'hc2 == req_index ? req_tag : tag_194; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1220 = 8'hc3 == req_index ? req_tag : tag_195; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1221 = 8'hc4 == req_index ? req_tag : tag_196; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1222 = 8'hc5 == req_index ? req_tag : tag_197; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1223 = 8'hc6 == req_index ? req_tag : tag_198; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1224 = 8'hc7 == req_index ? req_tag : tag_199; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1225 = 8'hc8 == req_index ? req_tag : tag_200; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1226 = 8'hc9 == req_index ? req_tag : tag_201; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1227 = 8'hca == req_index ? req_tag : tag_202; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1228 = 8'hcb == req_index ? req_tag : tag_203; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1229 = 8'hcc == req_index ? req_tag : tag_204; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1230 = 8'hcd == req_index ? req_tag : tag_205; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1231 = 8'hce == req_index ? req_tag : tag_206; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1232 = 8'hcf == req_index ? req_tag : tag_207; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1233 = 8'hd0 == req_index ? req_tag : tag_208; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1234 = 8'hd1 == req_index ? req_tag : tag_209; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1235 = 8'hd2 == req_index ? req_tag : tag_210; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1236 = 8'hd3 == req_index ? req_tag : tag_211; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1237 = 8'hd4 == req_index ? req_tag : tag_212; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1238 = 8'hd5 == req_index ? req_tag : tag_213; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1239 = 8'hd6 == req_index ? req_tag : tag_214; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1240 = 8'hd7 == req_index ? req_tag : tag_215; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1241 = 8'hd8 == req_index ? req_tag : tag_216; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1242 = 8'hd9 == req_index ? req_tag : tag_217; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1243 = 8'hda == req_index ? req_tag : tag_218; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1244 = 8'hdb == req_index ? req_tag : tag_219; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1245 = 8'hdc == req_index ? req_tag : tag_220; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1246 = 8'hdd == req_index ? req_tag : tag_221; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1247 = 8'hde == req_index ? req_tag : tag_222; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1248 = 8'hdf == req_index ? req_tag : tag_223; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1249 = 8'he0 == req_index ? req_tag : tag_224; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1250 = 8'he1 == req_index ? req_tag : tag_225; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1251 = 8'he2 == req_index ? req_tag : tag_226; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1252 = 8'he3 == req_index ? req_tag : tag_227; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1253 = 8'he4 == req_index ? req_tag : tag_228; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1254 = 8'he5 == req_index ? req_tag : tag_229; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1255 = 8'he6 == req_index ? req_tag : tag_230; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1256 = 8'he7 == req_index ? req_tag : tag_231; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1257 = 8'he8 == req_index ? req_tag : tag_232; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1258 = 8'he9 == req_index ? req_tag : tag_233; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1259 = 8'hea == req_index ? req_tag : tag_234; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1260 = 8'heb == req_index ? req_tag : tag_235; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1261 = 8'hec == req_index ? req_tag : tag_236; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1262 = 8'hed == req_index ? req_tag : tag_237; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1263 = 8'hee == req_index ? req_tag : tag_238; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1264 = 8'hef == req_index ? req_tag : tag_239; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1265 = 8'hf0 == req_index ? req_tag : tag_240; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1266 = 8'hf1 == req_index ? req_tag : tag_241; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1267 = 8'hf2 == req_index ? req_tag : tag_242; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1268 = 8'hf3 == req_index ? req_tag : tag_243; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1269 = 8'hf4 == req_index ? req_tag : tag_244; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1270 = 8'hf5 == req_index ? req_tag : tag_245; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1271 = 8'hf6 == req_index ? req_tag : tag_246; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1272 = 8'hf7 == req_index ? req_tag : tag_247; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1273 = 8'hf8 == req_index ? req_tag : tag_248; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1274 = 8'hf9 == req_index ? req_tag : tag_249; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1275 = 8'hfa == req_index ? req_tag : tag_250; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1276 = 8'hfb == req_index ? req_tag : tag_251; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1277 = 8'hfc == req_index ? req_tag : tag_252; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1278 = 8'hfd == req_index ? req_tag : tag_253; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1279 = 8'hfe == req_index ? req_tag : tag_254; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [19:0] _GEN_1280 = 8'hff == req_index ? req_tag : tag_255; // @[Dcache.scala 133:27 Dcache.scala 133:27 Dcache.scala 16:24]
  wire [3:0] _GEN_1281 = 8'h0 == req_index ? req_offset : offset_0; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1282 = 8'h1 == req_index ? req_offset : offset_1; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1283 = 8'h2 == req_index ? req_offset : offset_2; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1284 = 8'h3 == req_index ? req_offset : offset_3; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1285 = 8'h4 == req_index ? req_offset : offset_4; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1286 = 8'h5 == req_index ? req_offset : offset_5; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1287 = 8'h6 == req_index ? req_offset : offset_6; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1288 = 8'h7 == req_index ? req_offset : offset_7; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1289 = 8'h8 == req_index ? req_offset : offset_8; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1290 = 8'h9 == req_index ? req_offset : offset_9; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1291 = 8'ha == req_index ? req_offset : offset_10; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1292 = 8'hb == req_index ? req_offset : offset_11; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1293 = 8'hc == req_index ? req_offset : offset_12; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1294 = 8'hd == req_index ? req_offset : offset_13; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1295 = 8'he == req_index ? req_offset : offset_14; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1296 = 8'hf == req_index ? req_offset : offset_15; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1297 = 8'h10 == req_index ? req_offset : offset_16; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1298 = 8'h11 == req_index ? req_offset : offset_17; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1299 = 8'h12 == req_index ? req_offset : offset_18; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1300 = 8'h13 == req_index ? req_offset : offset_19; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1301 = 8'h14 == req_index ? req_offset : offset_20; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1302 = 8'h15 == req_index ? req_offset : offset_21; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1303 = 8'h16 == req_index ? req_offset : offset_22; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1304 = 8'h17 == req_index ? req_offset : offset_23; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1305 = 8'h18 == req_index ? req_offset : offset_24; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1306 = 8'h19 == req_index ? req_offset : offset_25; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1307 = 8'h1a == req_index ? req_offset : offset_26; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1308 = 8'h1b == req_index ? req_offset : offset_27; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1309 = 8'h1c == req_index ? req_offset : offset_28; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1310 = 8'h1d == req_index ? req_offset : offset_29; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1311 = 8'h1e == req_index ? req_offset : offset_30; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1312 = 8'h1f == req_index ? req_offset : offset_31; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1313 = 8'h20 == req_index ? req_offset : offset_32; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1314 = 8'h21 == req_index ? req_offset : offset_33; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1315 = 8'h22 == req_index ? req_offset : offset_34; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1316 = 8'h23 == req_index ? req_offset : offset_35; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1317 = 8'h24 == req_index ? req_offset : offset_36; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1318 = 8'h25 == req_index ? req_offset : offset_37; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1319 = 8'h26 == req_index ? req_offset : offset_38; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1320 = 8'h27 == req_index ? req_offset : offset_39; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1321 = 8'h28 == req_index ? req_offset : offset_40; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1322 = 8'h29 == req_index ? req_offset : offset_41; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1323 = 8'h2a == req_index ? req_offset : offset_42; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1324 = 8'h2b == req_index ? req_offset : offset_43; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1325 = 8'h2c == req_index ? req_offset : offset_44; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1326 = 8'h2d == req_index ? req_offset : offset_45; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1327 = 8'h2e == req_index ? req_offset : offset_46; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1328 = 8'h2f == req_index ? req_offset : offset_47; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1329 = 8'h30 == req_index ? req_offset : offset_48; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1330 = 8'h31 == req_index ? req_offset : offset_49; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1331 = 8'h32 == req_index ? req_offset : offset_50; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1332 = 8'h33 == req_index ? req_offset : offset_51; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1333 = 8'h34 == req_index ? req_offset : offset_52; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1334 = 8'h35 == req_index ? req_offset : offset_53; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1335 = 8'h36 == req_index ? req_offset : offset_54; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1336 = 8'h37 == req_index ? req_offset : offset_55; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1337 = 8'h38 == req_index ? req_offset : offset_56; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1338 = 8'h39 == req_index ? req_offset : offset_57; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1339 = 8'h3a == req_index ? req_offset : offset_58; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1340 = 8'h3b == req_index ? req_offset : offset_59; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1341 = 8'h3c == req_index ? req_offset : offset_60; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1342 = 8'h3d == req_index ? req_offset : offset_61; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1343 = 8'h3e == req_index ? req_offset : offset_62; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1344 = 8'h3f == req_index ? req_offset : offset_63; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1345 = 8'h40 == req_index ? req_offset : offset_64; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1346 = 8'h41 == req_index ? req_offset : offset_65; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1347 = 8'h42 == req_index ? req_offset : offset_66; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1348 = 8'h43 == req_index ? req_offset : offset_67; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1349 = 8'h44 == req_index ? req_offset : offset_68; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1350 = 8'h45 == req_index ? req_offset : offset_69; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1351 = 8'h46 == req_index ? req_offset : offset_70; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1352 = 8'h47 == req_index ? req_offset : offset_71; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1353 = 8'h48 == req_index ? req_offset : offset_72; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1354 = 8'h49 == req_index ? req_offset : offset_73; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1355 = 8'h4a == req_index ? req_offset : offset_74; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1356 = 8'h4b == req_index ? req_offset : offset_75; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1357 = 8'h4c == req_index ? req_offset : offset_76; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1358 = 8'h4d == req_index ? req_offset : offset_77; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1359 = 8'h4e == req_index ? req_offset : offset_78; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1360 = 8'h4f == req_index ? req_offset : offset_79; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1361 = 8'h50 == req_index ? req_offset : offset_80; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1362 = 8'h51 == req_index ? req_offset : offset_81; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1363 = 8'h52 == req_index ? req_offset : offset_82; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1364 = 8'h53 == req_index ? req_offset : offset_83; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1365 = 8'h54 == req_index ? req_offset : offset_84; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1366 = 8'h55 == req_index ? req_offset : offset_85; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1367 = 8'h56 == req_index ? req_offset : offset_86; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1368 = 8'h57 == req_index ? req_offset : offset_87; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1369 = 8'h58 == req_index ? req_offset : offset_88; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1370 = 8'h59 == req_index ? req_offset : offset_89; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1371 = 8'h5a == req_index ? req_offset : offset_90; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1372 = 8'h5b == req_index ? req_offset : offset_91; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1373 = 8'h5c == req_index ? req_offset : offset_92; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1374 = 8'h5d == req_index ? req_offset : offset_93; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1375 = 8'h5e == req_index ? req_offset : offset_94; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1376 = 8'h5f == req_index ? req_offset : offset_95; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1377 = 8'h60 == req_index ? req_offset : offset_96; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1378 = 8'h61 == req_index ? req_offset : offset_97; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1379 = 8'h62 == req_index ? req_offset : offset_98; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1380 = 8'h63 == req_index ? req_offset : offset_99; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1381 = 8'h64 == req_index ? req_offset : offset_100; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1382 = 8'h65 == req_index ? req_offset : offset_101; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1383 = 8'h66 == req_index ? req_offset : offset_102; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1384 = 8'h67 == req_index ? req_offset : offset_103; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1385 = 8'h68 == req_index ? req_offset : offset_104; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1386 = 8'h69 == req_index ? req_offset : offset_105; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1387 = 8'h6a == req_index ? req_offset : offset_106; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1388 = 8'h6b == req_index ? req_offset : offset_107; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1389 = 8'h6c == req_index ? req_offset : offset_108; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1390 = 8'h6d == req_index ? req_offset : offset_109; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1391 = 8'h6e == req_index ? req_offset : offset_110; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1392 = 8'h6f == req_index ? req_offset : offset_111; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1393 = 8'h70 == req_index ? req_offset : offset_112; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1394 = 8'h71 == req_index ? req_offset : offset_113; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1395 = 8'h72 == req_index ? req_offset : offset_114; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1396 = 8'h73 == req_index ? req_offset : offset_115; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1397 = 8'h74 == req_index ? req_offset : offset_116; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1398 = 8'h75 == req_index ? req_offset : offset_117; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1399 = 8'h76 == req_index ? req_offset : offset_118; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1400 = 8'h77 == req_index ? req_offset : offset_119; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1401 = 8'h78 == req_index ? req_offset : offset_120; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1402 = 8'h79 == req_index ? req_offset : offset_121; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1403 = 8'h7a == req_index ? req_offset : offset_122; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1404 = 8'h7b == req_index ? req_offset : offset_123; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1405 = 8'h7c == req_index ? req_offset : offset_124; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1406 = 8'h7d == req_index ? req_offset : offset_125; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1407 = 8'h7e == req_index ? req_offset : offset_126; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1408 = 8'h7f == req_index ? req_offset : offset_127; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1409 = 8'h80 == req_index ? req_offset : offset_128; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1410 = 8'h81 == req_index ? req_offset : offset_129; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1411 = 8'h82 == req_index ? req_offset : offset_130; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1412 = 8'h83 == req_index ? req_offset : offset_131; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1413 = 8'h84 == req_index ? req_offset : offset_132; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1414 = 8'h85 == req_index ? req_offset : offset_133; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1415 = 8'h86 == req_index ? req_offset : offset_134; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1416 = 8'h87 == req_index ? req_offset : offset_135; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1417 = 8'h88 == req_index ? req_offset : offset_136; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1418 = 8'h89 == req_index ? req_offset : offset_137; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1419 = 8'h8a == req_index ? req_offset : offset_138; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1420 = 8'h8b == req_index ? req_offset : offset_139; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1421 = 8'h8c == req_index ? req_offset : offset_140; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1422 = 8'h8d == req_index ? req_offset : offset_141; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1423 = 8'h8e == req_index ? req_offset : offset_142; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1424 = 8'h8f == req_index ? req_offset : offset_143; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1425 = 8'h90 == req_index ? req_offset : offset_144; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1426 = 8'h91 == req_index ? req_offset : offset_145; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1427 = 8'h92 == req_index ? req_offset : offset_146; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1428 = 8'h93 == req_index ? req_offset : offset_147; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1429 = 8'h94 == req_index ? req_offset : offset_148; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1430 = 8'h95 == req_index ? req_offset : offset_149; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1431 = 8'h96 == req_index ? req_offset : offset_150; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1432 = 8'h97 == req_index ? req_offset : offset_151; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1433 = 8'h98 == req_index ? req_offset : offset_152; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1434 = 8'h99 == req_index ? req_offset : offset_153; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1435 = 8'h9a == req_index ? req_offset : offset_154; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1436 = 8'h9b == req_index ? req_offset : offset_155; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1437 = 8'h9c == req_index ? req_offset : offset_156; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1438 = 8'h9d == req_index ? req_offset : offset_157; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1439 = 8'h9e == req_index ? req_offset : offset_158; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1440 = 8'h9f == req_index ? req_offset : offset_159; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1441 = 8'ha0 == req_index ? req_offset : offset_160; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1442 = 8'ha1 == req_index ? req_offset : offset_161; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1443 = 8'ha2 == req_index ? req_offset : offset_162; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1444 = 8'ha3 == req_index ? req_offset : offset_163; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1445 = 8'ha4 == req_index ? req_offset : offset_164; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1446 = 8'ha5 == req_index ? req_offset : offset_165; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1447 = 8'ha6 == req_index ? req_offset : offset_166; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1448 = 8'ha7 == req_index ? req_offset : offset_167; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1449 = 8'ha8 == req_index ? req_offset : offset_168; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1450 = 8'ha9 == req_index ? req_offset : offset_169; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1451 = 8'haa == req_index ? req_offset : offset_170; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1452 = 8'hab == req_index ? req_offset : offset_171; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1453 = 8'hac == req_index ? req_offset : offset_172; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1454 = 8'had == req_index ? req_offset : offset_173; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1455 = 8'hae == req_index ? req_offset : offset_174; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1456 = 8'haf == req_index ? req_offset : offset_175; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1457 = 8'hb0 == req_index ? req_offset : offset_176; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1458 = 8'hb1 == req_index ? req_offset : offset_177; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1459 = 8'hb2 == req_index ? req_offset : offset_178; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1460 = 8'hb3 == req_index ? req_offset : offset_179; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1461 = 8'hb4 == req_index ? req_offset : offset_180; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1462 = 8'hb5 == req_index ? req_offset : offset_181; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1463 = 8'hb6 == req_index ? req_offset : offset_182; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1464 = 8'hb7 == req_index ? req_offset : offset_183; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1465 = 8'hb8 == req_index ? req_offset : offset_184; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1466 = 8'hb9 == req_index ? req_offset : offset_185; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1467 = 8'hba == req_index ? req_offset : offset_186; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1468 = 8'hbb == req_index ? req_offset : offset_187; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1469 = 8'hbc == req_index ? req_offset : offset_188; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1470 = 8'hbd == req_index ? req_offset : offset_189; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1471 = 8'hbe == req_index ? req_offset : offset_190; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1472 = 8'hbf == req_index ? req_offset : offset_191; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1473 = 8'hc0 == req_index ? req_offset : offset_192; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1474 = 8'hc1 == req_index ? req_offset : offset_193; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1475 = 8'hc2 == req_index ? req_offset : offset_194; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1476 = 8'hc3 == req_index ? req_offset : offset_195; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1477 = 8'hc4 == req_index ? req_offset : offset_196; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1478 = 8'hc5 == req_index ? req_offset : offset_197; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1479 = 8'hc6 == req_index ? req_offset : offset_198; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1480 = 8'hc7 == req_index ? req_offset : offset_199; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1481 = 8'hc8 == req_index ? req_offset : offset_200; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1482 = 8'hc9 == req_index ? req_offset : offset_201; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1483 = 8'hca == req_index ? req_offset : offset_202; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1484 = 8'hcb == req_index ? req_offset : offset_203; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1485 = 8'hcc == req_index ? req_offset : offset_204; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1486 = 8'hcd == req_index ? req_offset : offset_205; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1487 = 8'hce == req_index ? req_offset : offset_206; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1488 = 8'hcf == req_index ? req_offset : offset_207; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1489 = 8'hd0 == req_index ? req_offset : offset_208; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1490 = 8'hd1 == req_index ? req_offset : offset_209; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1491 = 8'hd2 == req_index ? req_offset : offset_210; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1492 = 8'hd3 == req_index ? req_offset : offset_211; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1493 = 8'hd4 == req_index ? req_offset : offset_212; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1494 = 8'hd5 == req_index ? req_offset : offset_213; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1495 = 8'hd6 == req_index ? req_offset : offset_214; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1496 = 8'hd7 == req_index ? req_offset : offset_215; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1497 = 8'hd8 == req_index ? req_offset : offset_216; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1498 = 8'hd9 == req_index ? req_offset : offset_217; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1499 = 8'hda == req_index ? req_offset : offset_218; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1500 = 8'hdb == req_index ? req_offset : offset_219; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1501 = 8'hdc == req_index ? req_offset : offset_220; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1502 = 8'hdd == req_index ? req_offset : offset_221; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1503 = 8'hde == req_index ? req_offset : offset_222; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1504 = 8'hdf == req_index ? req_offset : offset_223; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1505 = 8'he0 == req_index ? req_offset : offset_224; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1506 = 8'he1 == req_index ? req_offset : offset_225; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1507 = 8'he2 == req_index ? req_offset : offset_226; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1508 = 8'he3 == req_index ? req_offset : offset_227; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1509 = 8'he4 == req_index ? req_offset : offset_228; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1510 = 8'he5 == req_index ? req_offset : offset_229; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1511 = 8'he6 == req_index ? req_offset : offset_230; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1512 = 8'he7 == req_index ? req_offset : offset_231; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1513 = 8'he8 == req_index ? req_offset : offset_232; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1514 = 8'he9 == req_index ? req_offset : offset_233; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1515 = 8'hea == req_index ? req_offset : offset_234; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1516 = 8'heb == req_index ? req_offset : offset_235; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1517 = 8'hec == req_index ? req_offset : offset_236; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1518 = 8'hed == req_index ? req_offset : offset_237; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1519 = 8'hee == req_index ? req_offset : offset_238; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1520 = 8'hef == req_index ? req_offset : offset_239; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1521 = 8'hf0 == req_index ? req_offset : offset_240; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1522 = 8'hf1 == req_index ? req_offset : offset_241; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1523 = 8'hf2 == req_index ? req_offset : offset_242; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1524 = 8'hf3 == req_index ? req_offset : offset_243; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1525 = 8'hf4 == req_index ? req_offset : offset_244; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1526 = 8'hf5 == req_index ? req_offset : offset_245; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1527 = 8'hf6 == req_index ? req_offset : offset_246; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1528 = 8'hf7 == req_index ? req_offset : offset_247; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1529 = 8'hf8 == req_index ? req_offset : offset_248; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1530 = 8'hf9 == req_index ? req_offset : offset_249; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1531 = 8'hfa == req_index ? req_offset : offset_250; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1532 = 8'hfb == req_index ? req_offset : offset_251; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1533 = 8'hfc == req_index ? req_offset : offset_252; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1534 = 8'hfd == req_index ? req_offset : offset_253; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1535 = 8'hfe == req_index ? req_offset : offset_254; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [3:0] _GEN_1536 = 8'hff == req_index ? req_offset : offset_255; // @[Dcache.scala 134:27 Dcache.scala 134:27 Dcache.scala 19:24]
  wire [127:0] _cache_wdata_T_1 = {valid_wdata,64'h0}; // @[Cat.scala 30:58]
  wire [127:0] _cache_wdata_T_2 = {64'h0,valid_wdata}; // @[Cat.scala 30:58]
  wire [127:0] _cache_wdata_T_3 = req_offset[3] ? _cache_wdata_T_1 : _cache_wdata_T_2; // @[Dcache.scala 137:33]
  wire [127:0] _cache_strb_T_1 = {valid_strb,64'h0}; // @[Cat.scala 30:58]
  wire [127:0] _cache_strb_T_2 = {64'h0,valid_strb}; // @[Cat.scala 30:58]
  wire [127:0] _cache_strb_T_3 = req_offset[3] ? _cache_strb_T_1 : _cache_strb_T_2; // @[Dcache.scala 138:33]
  wire  _GEN_1537 = 8'h0 == req_index ? io_dmem_data_req : dirty_0; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1538 = 8'h1 == req_index ? io_dmem_data_req : dirty_1; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1539 = 8'h2 == req_index ? io_dmem_data_req : dirty_2; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1540 = 8'h3 == req_index ? io_dmem_data_req : dirty_3; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1541 = 8'h4 == req_index ? io_dmem_data_req : dirty_4; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1542 = 8'h5 == req_index ? io_dmem_data_req : dirty_5; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1543 = 8'h6 == req_index ? io_dmem_data_req : dirty_6; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1544 = 8'h7 == req_index ? io_dmem_data_req : dirty_7; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1545 = 8'h8 == req_index ? io_dmem_data_req : dirty_8; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1546 = 8'h9 == req_index ? io_dmem_data_req : dirty_9; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1547 = 8'ha == req_index ? io_dmem_data_req : dirty_10; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1548 = 8'hb == req_index ? io_dmem_data_req : dirty_11; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1549 = 8'hc == req_index ? io_dmem_data_req : dirty_12; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1550 = 8'hd == req_index ? io_dmem_data_req : dirty_13; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1551 = 8'he == req_index ? io_dmem_data_req : dirty_14; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1552 = 8'hf == req_index ? io_dmem_data_req : dirty_15; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1553 = 8'h10 == req_index ? io_dmem_data_req : dirty_16; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1554 = 8'h11 == req_index ? io_dmem_data_req : dirty_17; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1555 = 8'h12 == req_index ? io_dmem_data_req : dirty_18; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1556 = 8'h13 == req_index ? io_dmem_data_req : dirty_19; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1557 = 8'h14 == req_index ? io_dmem_data_req : dirty_20; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1558 = 8'h15 == req_index ? io_dmem_data_req : dirty_21; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1559 = 8'h16 == req_index ? io_dmem_data_req : dirty_22; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1560 = 8'h17 == req_index ? io_dmem_data_req : dirty_23; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1561 = 8'h18 == req_index ? io_dmem_data_req : dirty_24; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1562 = 8'h19 == req_index ? io_dmem_data_req : dirty_25; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1563 = 8'h1a == req_index ? io_dmem_data_req : dirty_26; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1564 = 8'h1b == req_index ? io_dmem_data_req : dirty_27; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1565 = 8'h1c == req_index ? io_dmem_data_req : dirty_28; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1566 = 8'h1d == req_index ? io_dmem_data_req : dirty_29; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1567 = 8'h1e == req_index ? io_dmem_data_req : dirty_30; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1568 = 8'h1f == req_index ? io_dmem_data_req : dirty_31; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1569 = 8'h20 == req_index ? io_dmem_data_req : dirty_32; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1570 = 8'h21 == req_index ? io_dmem_data_req : dirty_33; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1571 = 8'h22 == req_index ? io_dmem_data_req : dirty_34; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1572 = 8'h23 == req_index ? io_dmem_data_req : dirty_35; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1573 = 8'h24 == req_index ? io_dmem_data_req : dirty_36; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1574 = 8'h25 == req_index ? io_dmem_data_req : dirty_37; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1575 = 8'h26 == req_index ? io_dmem_data_req : dirty_38; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1576 = 8'h27 == req_index ? io_dmem_data_req : dirty_39; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1577 = 8'h28 == req_index ? io_dmem_data_req : dirty_40; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1578 = 8'h29 == req_index ? io_dmem_data_req : dirty_41; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1579 = 8'h2a == req_index ? io_dmem_data_req : dirty_42; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1580 = 8'h2b == req_index ? io_dmem_data_req : dirty_43; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1581 = 8'h2c == req_index ? io_dmem_data_req : dirty_44; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1582 = 8'h2d == req_index ? io_dmem_data_req : dirty_45; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1583 = 8'h2e == req_index ? io_dmem_data_req : dirty_46; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1584 = 8'h2f == req_index ? io_dmem_data_req : dirty_47; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1585 = 8'h30 == req_index ? io_dmem_data_req : dirty_48; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1586 = 8'h31 == req_index ? io_dmem_data_req : dirty_49; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1587 = 8'h32 == req_index ? io_dmem_data_req : dirty_50; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1588 = 8'h33 == req_index ? io_dmem_data_req : dirty_51; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1589 = 8'h34 == req_index ? io_dmem_data_req : dirty_52; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1590 = 8'h35 == req_index ? io_dmem_data_req : dirty_53; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1591 = 8'h36 == req_index ? io_dmem_data_req : dirty_54; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1592 = 8'h37 == req_index ? io_dmem_data_req : dirty_55; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1593 = 8'h38 == req_index ? io_dmem_data_req : dirty_56; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1594 = 8'h39 == req_index ? io_dmem_data_req : dirty_57; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1595 = 8'h3a == req_index ? io_dmem_data_req : dirty_58; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1596 = 8'h3b == req_index ? io_dmem_data_req : dirty_59; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1597 = 8'h3c == req_index ? io_dmem_data_req : dirty_60; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1598 = 8'h3d == req_index ? io_dmem_data_req : dirty_61; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1599 = 8'h3e == req_index ? io_dmem_data_req : dirty_62; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1600 = 8'h3f == req_index ? io_dmem_data_req : dirty_63; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1601 = 8'h40 == req_index ? io_dmem_data_req : dirty_64; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1602 = 8'h41 == req_index ? io_dmem_data_req : dirty_65; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1603 = 8'h42 == req_index ? io_dmem_data_req : dirty_66; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1604 = 8'h43 == req_index ? io_dmem_data_req : dirty_67; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1605 = 8'h44 == req_index ? io_dmem_data_req : dirty_68; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1606 = 8'h45 == req_index ? io_dmem_data_req : dirty_69; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1607 = 8'h46 == req_index ? io_dmem_data_req : dirty_70; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1608 = 8'h47 == req_index ? io_dmem_data_req : dirty_71; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1609 = 8'h48 == req_index ? io_dmem_data_req : dirty_72; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1610 = 8'h49 == req_index ? io_dmem_data_req : dirty_73; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1611 = 8'h4a == req_index ? io_dmem_data_req : dirty_74; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1612 = 8'h4b == req_index ? io_dmem_data_req : dirty_75; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1613 = 8'h4c == req_index ? io_dmem_data_req : dirty_76; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1614 = 8'h4d == req_index ? io_dmem_data_req : dirty_77; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1615 = 8'h4e == req_index ? io_dmem_data_req : dirty_78; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1616 = 8'h4f == req_index ? io_dmem_data_req : dirty_79; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1617 = 8'h50 == req_index ? io_dmem_data_req : dirty_80; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1618 = 8'h51 == req_index ? io_dmem_data_req : dirty_81; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1619 = 8'h52 == req_index ? io_dmem_data_req : dirty_82; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1620 = 8'h53 == req_index ? io_dmem_data_req : dirty_83; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1621 = 8'h54 == req_index ? io_dmem_data_req : dirty_84; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1622 = 8'h55 == req_index ? io_dmem_data_req : dirty_85; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1623 = 8'h56 == req_index ? io_dmem_data_req : dirty_86; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1624 = 8'h57 == req_index ? io_dmem_data_req : dirty_87; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1625 = 8'h58 == req_index ? io_dmem_data_req : dirty_88; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1626 = 8'h59 == req_index ? io_dmem_data_req : dirty_89; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1627 = 8'h5a == req_index ? io_dmem_data_req : dirty_90; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1628 = 8'h5b == req_index ? io_dmem_data_req : dirty_91; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1629 = 8'h5c == req_index ? io_dmem_data_req : dirty_92; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1630 = 8'h5d == req_index ? io_dmem_data_req : dirty_93; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1631 = 8'h5e == req_index ? io_dmem_data_req : dirty_94; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1632 = 8'h5f == req_index ? io_dmem_data_req : dirty_95; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1633 = 8'h60 == req_index ? io_dmem_data_req : dirty_96; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1634 = 8'h61 == req_index ? io_dmem_data_req : dirty_97; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1635 = 8'h62 == req_index ? io_dmem_data_req : dirty_98; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1636 = 8'h63 == req_index ? io_dmem_data_req : dirty_99; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1637 = 8'h64 == req_index ? io_dmem_data_req : dirty_100; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1638 = 8'h65 == req_index ? io_dmem_data_req : dirty_101; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1639 = 8'h66 == req_index ? io_dmem_data_req : dirty_102; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1640 = 8'h67 == req_index ? io_dmem_data_req : dirty_103; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1641 = 8'h68 == req_index ? io_dmem_data_req : dirty_104; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1642 = 8'h69 == req_index ? io_dmem_data_req : dirty_105; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1643 = 8'h6a == req_index ? io_dmem_data_req : dirty_106; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1644 = 8'h6b == req_index ? io_dmem_data_req : dirty_107; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1645 = 8'h6c == req_index ? io_dmem_data_req : dirty_108; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1646 = 8'h6d == req_index ? io_dmem_data_req : dirty_109; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1647 = 8'h6e == req_index ? io_dmem_data_req : dirty_110; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1648 = 8'h6f == req_index ? io_dmem_data_req : dirty_111; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1649 = 8'h70 == req_index ? io_dmem_data_req : dirty_112; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1650 = 8'h71 == req_index ? io_dmem_data_req : dirty_113; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1651 = 8'h72 == req_index ? io_dmem_data_req : dirty_114; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1652 = 8'h73 == req_index ? io_dmem_data_req : dirty_115; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1653 = 8'h74 == req_index ? io_dmem_data_req : dirty_116; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1654 = 8'h75 == req_index ? io_dmem_data_req : dirty_117; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1655 = 8'h76 == req_index ? io_dmem_data_req : dirty_118; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1656 = 8'h77 == req_index ? io_dmem_data_req : dirty_119; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1657 = 8'h78 == req_index ? io_dmem_data_req : dirty_120; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1658 = 8'h79 == req_index ? io_dmem_data_req : dirty_121; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1659 = 8'h7a == req_index ? io_dmem_data_req : dirty_122; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1660 = 8'h7b == req_index ? io_dmem_data_req : dirty_123; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1661 = 8'h7c == req_index ? io_dmem_data_req : dirty_124; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1662 = 8'h7d == req_index ? io_dmem_data_req : dirty_125; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1663 = 8'h7e == req_index ? io_dmem_data_req : dirty_126; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1664 = 8'h7f == req_index ? io_dmem_data_req : dirty_127; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1665 = 8'h80 == req_index ? io_dmem_data_req : dirty_128; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1666 = 8'h81 == req_index ? io_dmem_data_req : dirty_129; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1667 = 8'h82 == req_index ? io_dmem_data_req : dirty_130; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1668 = 8'h83 == req_index ? io_dmem_data_req : dirty_131; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1669 = 8'h84 == req_index ? io_dmem_data_req : dirty_132; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1670 = 8'h85 == req_index ? io_dmem_data_req : dirty_133; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1671 = 8'h86 == req_index ? io_dmem_data_req : dirty_134; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1672 = 8'h87 == req_index ? io_dmem_data_req : dirty_135; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1673 = 8'h88 == req_index ? io_dmem_data_req : dirty_136; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1674 = 8'h89 == req_index ? io_dmem_data_req : dirty_137; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1675 = 8'h8a == req_index ? io_dmem_data_req : dirty_138; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1676 = 8'h8b == req_index ? io_dmem_data_req : dirty_139; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1677 = 8'h8c == req_index ? io_dmem_data_req : dirty_140; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1678 = 8'h8d == req_index ? io_dmem_data_req : dirty_141; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1679 = 8'h8e == req_index ? io_dmem_data_req : dirty_142; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1680 = 8'h8f == req_index ? io_dmem_data_req : dirty_143; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1681 = 8'h90 == req_index ? io_dmem_data_req : dirty_144; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1682 = 8'h91 == req_index ? io_dmem_data_req : dirty_145; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1683 = 8'h92 == req_index ? io_dmem_data_req : dirty_146; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1684 = 8'h93 == req_index ? io_dmem_data_req : dirty_147; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1685 = 8'h94 == req_index ? io_dmem_data_req : dirty_148; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1686 = 8'h95 == req_index ? io_dmem_data_req : dirty_149; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1687 = 8'h96 == req_index ? io_dmem_data_req : dirty_150; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1688 = 8'h97 == req_index ? io_dmem_data_req : dirty_151; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1689 = 8'h98 == req_index ? io_dmem_data_req : dirty_152; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1690 = 8'h99 == req_index ? io_dmem_data_req : dirty_153; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1691 = 8'h9a == req_index ? io_dmem_data_req : dirty_154; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1692 = 8'h9b == req_index ? io_dmem_data_req : dirty_155; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1693 = 8'h9c == req_index ? io_dmem_data_req : dirty_156; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1694 = 8'h9d == req_index ? io_dmem_data_req : dirty_157; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1695 = 8'h9e == req_index ? io_dmem_data_req : dirty_158; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1696 = 8'h9f == req_index ? io_dmem_data_req : dirty_159; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1697 = 8'ha0 == req_index ? io_dmem_data_req : dirty_160; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1698 = 8'ha1 == req_index ? io_dmem_data_req : dirty_161; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1699 = 8'ha2 == req_index ? io_dmem_data_req : dirty_162; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1700 = 8'ha3 == req_index ? io_dmem_data_req : dirty_163; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1701 = 8'ha4 == req_index ? io_dmem_data_req : dirty_164; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1702 = 8'ha5 == req_index ? io_dmem_data_req : dirty_165; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1703 = 8'ha6 == req_index ? io_dmem_data_req : dirty_166; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1704 = 8'ha7 == req_index ? io_dmem_data_req : dirty_167; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1705 = 8'ha8 == req_index ? io_dmem_data_req : dirty_168; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1706 = 8'ha9 == req_index ? io_dmem_data_req : dirty_169; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1707 = 8'haa == req_index ? io_dmem_data_req : dirty_170; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1708 = 8'hab == req_index ? io_dmem_data_req : dirty_171; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1709 = 8'hac == req_index ? io_dmem_data_req : dirty_172; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1710 = 8'had == req_index ? io_dmem_data_req : dirty_173; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1711 = 8'hae == req_index ? io_dmem_data_req : dirty_174; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1712 = 8'haf == req_index ? io_dmem_data_req : dirty_175; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1713 = 8'hb0 == req_index ? io_dmem_data_req : dirty_176; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1714 = 8'hb1 == req_index ? io_dmem_data_req : dirty_177; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1715 = 8'hb2 == req_index ? io_dmem_data_req : dirty_178; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1716 = 8'hb3 == req_index ? io_dmem_data_req : dirty_179; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1717 = 8'hb4 == req_index ? io_dmem_data_req : dirty_180; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1718 = 8'hb5 == req_index ? io_dmem_data_req : dirty_181; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1719 = 8'hb6 == req_index ? io_dmem_data_req : dirty_182; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1720 = 8'hb7 == req_index ? io_dmem_data_req : dirty_183; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1721 = 8'hb8 == req_index ? io_dmem_data_req : dirty_184; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1722 = 8'hb9 == req_index ? io_dmem_data_req : dirty_185; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1723 = 8'hba == req_index ? io_dmem_data_req : dirty_186; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1724 = 8'hbb == req_index ? io_dmem_data_req : dirty_187; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1725 = 8'hbc == req_index ? io_dmem_data_req : dirty_188; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1726 = 8'hbd == req_index ? io_dmem_data_req : dirty_189; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1727 = 8'hbe == req_index ? io_dmem_data_req : dirty_190; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1728 = 8'hbf == req_index ? io_dmem_data_req : dirty_191; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1729 = 8'hc0 == req_index ? io_dmem_data_req : dirty_192; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1730 = 8'hc1 == req_index ? io_dmem_data_req : dirty_193; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1731 = 8'hc2 == req_index ? io_dmem_data_req : dirty_194; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1732 = 8'hc3 == req_index ? io_dmem_data_req : dirty_195; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1733 = 8'hc4 == req_index ? io_dmem_data_req : dirty_196; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1734 = 8'hc5 == req_index ? io_dmem_data_req : dirty_197; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1735 = 8'hc6 == req_index ? io_dmem_data_req : dirty_198; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1736 = 8'hc7 == req_index ? io_dmem_data_req : dirty_199; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1737 = 8'hc8 == req_index ? io_dmem_data_req : dirty_200; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1738 = 8'hc9 == req_index ? io_dmem_data_req : dirty_201; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1739 = 8'hca == req_index ? io_dmem_data_req : dirty_202; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1740 = 8'hcb == req_index ? io_dmem_data_req : dirty_203; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1741 = 8'hcc == req_index ? io_dmem_data_req : dirty_204; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1742 = 8'hcd == req_index ? io_dmem_data_req : dirty_205; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1743 = 8'hce == req_index ? io_dmem_data_req : dirty_206; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1744 = 8'hcf == req_index ? io_dmem_data_req : dirty_207; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1745 = 8'hd0 == req_index ? io_dmem_data_req : dirty_208; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1746 = 8'hd1 == req_index ? io_dmem_data_req : dirty_209; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1747 = 8'hd2 == req_index ? io_dmem_data_req : dirty_210; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1748 = 8'hd3 == req_index ? io_dmem_data_req : dirty_211; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1749 = 8'hd4 == req_index ? io_dmem_data_req : dirty_212; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1750 = 8'hd5 == req_index ? io_dmem_data_req : dirty_213; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1751 = 8'hd6 == req_index ? io_dmem_data_req : dirty_214; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1752 = 8'hd7 == req_index ? io_dmem_data_req : dirty_215; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1753 = 8'hd8 == req_index ? io_dmem_data_req : dirty_216; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1754 = 8'hd9 == req_index ? io_dmem_data_req : dirty_217; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1755 = 8'hda == req_index ? io_dmem_data_req : dirty_218; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1756 = 8'hdb == req_index ? io_dmem_data_req : dirty_219; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1757 = 8'hdc == req_index ? io_dmem_data_req : dirty_220; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1758 = 8'hdd == req_index ? io_dmem_data_req : dirty_221; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1759 = 8'hde == req_index ? io_dmem_data_req : dirty_222; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1760 = 8'hdf == req_index ? io_dmem_data_req : dirty_223; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1761 = 8'he0 == req_index ? io_dmem_data_req : dirty_224; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1762 = 8'he1 == req_index ? io_dmem_data_req : dirty_225; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1763 = 8'he2 == req_index ? io_dmem_data_req : dirty_226; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1764 = 8'he3 == req_index ? io_dmem_data_req : dirty_227; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1765 = 8'he4 == req_index ? io_dmem_data_req : dirty_228; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1766 = 8'he5 == req_index ? io_dmem_data_req : dirty_229; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1767 = 8'he6 == req_index ? io_dmem_data_req : dirty_230; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1768 = 8'he7 == req_index ? io_dmem_data_req : dirty_231; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1769 = 8'he8 == req_index ? io_dmem_data_req : dirty_232; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1770 = 8'he9 == req_index ? io_dmem_data_req : dirty_233; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1771 = 8'hea == req_index ? io_dmem_data_req : dirty_234; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1772 = 8'heb == req_index ? io_dmem_data_req : dirty_235; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1773 = 8'hec == req_index ? io_dmem_data_req : dirty_236; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1774 = 8'hed == req_index ? io_dmem_data_req : dirty_237; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1775 = 8'hee == req_index ? io_dmem_data_req : dirty_238; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1776 = 8'hef == req_index ? io_dmem_data_req : dirty_239; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1777 = 8'hf0 == req_index ? io_dmem_data_req : dirty_240; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1778 = 8'hf1 == req_index ? io_dmem_data_req : dirty_241; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1779 = 8'hf2 == req_index ? io_dmem_data_req : dirty_242; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1780 = 8'hf3 == req_index ? io_dmem_data_req : dirty_243; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1781 = 8'hf4 == req_index ? io_dmem_data_req : dirty_244; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1782 = 8'hf5 == req_index ? io_dmem_data_req : dirty_245; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1783 = 8'hf6 == req_index ? io_dmem_data_req : dirty_246; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1784 = 8'hf7 == req_index ? io_dmem_data_req : dirty_247; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1785 = 8'hf8 == req_index ? io_dmem_data_req : dirty_248; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1786 = 8'hf9 == req_index ? io_dmem_data_req : dirty_249; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1787 = 8'hfa == req_index ? io_dmem_data_req : dirty_250; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1788 = 8'hfb == req_index ? io_dmem_data_req : dirty_251; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1789 = 8'hfc == req_index ? io_dmem_data_req : dirty_252; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1790 = 8'hfd == req_index ? io_dmem_data_req : dirty_253; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1791 = 8'hfe == req_index ? io_dmem_data_req : dirty_254; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1792 = 8'hff == req_index ? io_dmem_data_req : dirty_255; // @[Dcache.scala 140:28 Dcache.scala 140:28 Dcache.scala 18:24]
  wire  _GEN_1793 = ~_GEN_767 ? _GEN_1537 : dirty_0; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1794 = ~_GEN_767 ? _GEN_1538 : dirty_1; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1795 = ~_GEN_767 ? _GEN_1539 : dirty_2; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1796 = ~_GEN_767 ? _GEN_1540 : dirty_3; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1797 = ~_GEN_767 ? _GEN_1541 : dirty_4; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1798 = ~_GEN_767 ? _GEN_1542 : dirty_5; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1799 = ~_GEN_767 ? _GEN_1543 : dirty_6; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1800 = ~_GEN_767 ? _GEN_1544 : dirty_7; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1801 = ~_GEN_767 ? _GEN_1545 : dirty_8; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1802 = ~_GEN_767 ? _GEN_1546 : dirty_9; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1803 = ~_GEN_767 ? _GEN_1547 : dirty_10; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1804 = ~_GEN_767 ? _GEN_1548 : dirty_11; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1805 = ~_GEN_767 ? _GEN_1549 : dirty_12; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1806 = ~_GEN_767 ? _GEN_1550 : dirty_13; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1807 = ~_GEN_767 ? _GEN_1551 : dirty_14; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1808 = ~_GEN_767 ? _GEN_1552 : dirty_15; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1809 = ~_GEN_767 ? _GEN_1553 : dirty_16; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1810 = ~_GEN_767 ? _GEN_1554 : dirty_17; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1811 = ~_GEN_767 ? _GEN_1555 : dirty_18; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1812 = ~_GEN_767 ? _GEN_1556 : dirty_19; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1813 = ~_GEN_767 ? _GEN_1557 : dirty_20; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1814 = ~_GEN_767 ? _GEN_1558 : dirty_21; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1815 = ~_GEN_767 ? _GEN_1559 : dirty_22; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1816 = ~_GEN_767 ? _GEN_1560 : dirty_23; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1817 = ~_GEN_767 ? _GEN_1561 : dirty_24; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1818 = ~_GEN_767 ? _GEN_1562 : dirty_25; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1819 = ~_GEN_767 ? _GEN_1563 : dirty_26; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1820 = ~_GEN_767 ? _GEN_1564 : dirty_27; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1821 = ~_GEN_767 ? _GEN_1565 : dirty_28; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1822 = ~_GEN_767 ? _GEN_1566 : dirty_29; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1823 = ~_GEN_767 ? _GEN_1567 : dirty_30; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1824 = ~_GEN_767 ? _GEN_1568 : dirty_31; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1825 = ~_GEN_767 ? _GEN_1569 : dirty_32; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1826 = ~_GEN_767 ? _GEN_1570 : dirty_33; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1827 = ~_GEN_767 ? _GEN_1571 : dirty_34; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1828 = ~_GEN_767 ? _GEN_1572 : dirty_35; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1829 = ~_GEN_767 ? _GEN_1573 : dirty_36; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1830 = ~_GEN_767 ? _GEN_1574 : dirty_37; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1831 = ~_GEN_767 ? _GEN_1575 : dirty_38; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1832 = ~_GEN_767 ? _GEN_1576 : dirty_39; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1833 = ~_GEN_767 ? _GEN_1577 : dirty_40; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1834 = ~_GEN_767 ? _GEN_1578 : dirty_41; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1835 = ~_GEN_767 ? _GEN_1579 : dirty_42; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1836 = ~_GEN_767 ? _GEN_1580 : dirty_43; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1837 = ~_GEN_767 ? _GEN_1581 : dirty_44; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1838 = ~_GEN_767 ? _GEN_1582 : dirty_45; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1839 = ~_GEN_767 ? _GEN_1583 : dirty_46; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1840 = ~_GEN_767 ? _GEN_1584 : dirty_47; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1841 = ~_GEN_767 ? _GEN_1585 : dirty_48; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1842 = ~_GEN_767 ? _GEN_1586 : dirty_49; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1843 = ~_GEN_767 ? _GEN_1587 : dirty_50; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1844 = ~_GEN_767 ? _GEN_1588 : dirty_51; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1845 = ~_GEN_767 ? _GEN_1589 : dirty_52; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1846 = ~_GEN_767 ? _GEN_1590 : dirty_53; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1847 = ~_GEN_767 ? _GEN_1591 : dirty_54; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1848 = ~_GEN_767 ? _GEN_1592 : dirty_55; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1849 = ~_GEN_767 ? _GEN_1593 : dirty_56; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1850 = ~_GEN_767 ? _GEN_1594 : dirty_57; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1851 = ~_GEN_767 ? _GEN_1595 : dirty_58; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1852 = ~_GEN_767 ? _GEN_1596 : dirty_59; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1853 = ~_GEN_767 ? _GEN_1597 : dirty_60; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1854 = ~_GEN_767 ? _GEN_1598 : dirty_61; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1855 = ~_GEN_767 ? _GEN_1599 : dirty_62; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1856 = ~_GEN_767 ? _GEN_1600 : dirty_63; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1857 = ~_GEN_767 ? _GEN_1601 : dirty_64; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1858 = ~_GEN_767 ? _GEN_1602 : dirty_65; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1859 = ~_GEN_767 ? _GEN_1603 : dirty_66; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1860 = ~_GEN_767 ? _GEN_1604 : dirty_67; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1861 = ~_GEN_767 ? _GEN_1605 : dirty_68; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1862 = ~_GEN_767 ? _GEN_1606 : dirty_69; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1863 = ~_GEN_767 ? _GEN_1607 : dirty_70; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1864 = ~_GEN_767 ? _GEN_1608 : dirty_71; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1865 = ~_GEN_767 ? _GEN_1609 : dirty_72; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1866 = ~_GEN_767 ? _GEN_1610 : dirty_73; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1867 = ~_GEN_767 ? _GEN_1611 : dirty_74; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1868 = ~_GEN_767 ? _GEN_1612 : dirty_75; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1869 = ~_GEN_767 ? _GEN_1613 : dirty_76; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1870 = ~_GEN_767 ? _GEN_1614 : dirty_77; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1871 = ~_GEN_767 ? _GEN_1615 : dirty_78; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1872 = ~_GEN_767 ? _GEN_1616 : dirty_79; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1873 = ~_GEN_767 ? _GEN_1617 : dirty_80; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1874 = ~_GEN_767 ? _GEN_1618 : dirty_81; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1875 = ~_GEN_767 ? _GEN_1619 : dirty_82; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1876 = ~_GEN_767 ? _GEN_1620 : dirty_83; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1877 = ~_GEN_767 ? _GEN_1621 : dirty_84; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1878 = ~_GEN_767 ? _GEN_1622 : dirty_85; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1879 = ~_GEN_767 ? _GEN_1623 : dirty_86; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1880 = ~_GEN_767 ? _GEN_1624 : dirty_87; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1881 = ~_GEN_767 ? _GEN_1625 : dirty_88; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1882 = ~_GEN_767 ? _GEN_1626 : dirty_89; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1883 = ~_GEN_767 ? _GEN_1627 : dirty_90; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1884 = ~_GEN_767 ? _GEN_1628 : dirty_91; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1885 = ~_GEN_767 ? _GEN_1629 : dirty_92; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1886 = ~_GEN_767 ? _GEN_1630 : dirty_93; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1887 = ~_GEN_767 ? _GEN_1631 : dirty_94; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1888 = ~_GEN_767 ? _GEN_1632 : dirty_95; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1889 = ~_GEN_767 ? _GEN_1633 : dirty_96; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1890 = ~_GEN_767 ? _GEN_1634 : dirty_97; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1891 = ~_GEN_767 ? _GEN_1635 : dirty_98; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1892 = ~_GEN_767 ? _GEN_1636 : dirty_99; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1893 = ~_GEN_767 ? _GEN_1637 : dirty_100; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1894 = ~_GEN_767 ? _GEN_1638 : dirty_101; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1895 = ~_GEN_767 ? _GEN_1639 : dirty_102; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1896 = ~_GEN_767 ? _GEN_1640 : dirty_103; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1897 = ~_GEN_767 ? _GEN_1641 : dirty_104; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1898 = ~_GEN_767 ? _GEN_1642 : dirty_105; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1899 = ~_GEN_767 ? _GEN_1643 : dirty_106; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1900 = ~_GEN_767 ? _GEN_1644 : dirty_107; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1901 = ~_GEN_767 ? _GEN_1645 : dirty_108; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1902 = ~_GEN_767 ? _GEN_1646 : dirty_109; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1903 = ~_GEN_767 ? _GEN_1647 : dirty_110; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1904 = ~_GEN_767 ? _GEN_1648 : dirty_111; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1905 = ~_GEN_767 ? _GEN_1649 : dirty_112; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1906 = ~_GEN_767 ? _GEN_1650 : dirty_113; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1907 = ~_GEN_767 ? _GEN_1651 : dirty_114; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1908 = ~_GEN_767 ? _GEN_1652 : dirty_115; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1909 = ~_GEN_767 ? _GEN_1653 : dirty_116; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1910 = ~_GEN_767 ? _GEN_1654 : dirty_117; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1911 = ~_GEN_767 ? _GEN_1655 : dirty_118; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1912 = ~_GEN_767 ? _GEN_1656 : dirty_119; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1913 = ~_GEN_767 ? _GEN_1657 : dirty_120; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1914 = ~_GEN_767 ? _GEN_1658 : dirty_121; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1915 = ~_GEN_767 ? _GEN_1659 : dirty_122; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1916 = ~_GEN_767 ? _GEN_1660 : dirty_123; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1917 = ~_GEN_767 ? _GEN_1661 : dirty_124; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1918 = ~_GEN_767 ? _GEN_1662 : dirty_125; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1919 = ~_GEN_767 ? _GEN_1663 : dirty_126; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1920 = ~_GEN_767 ? _GEN_1664 : dirty_127; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1921 = ~_GEN_767 ? _GEN_1665 : dirty_128; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1922 = ~_GEN_767 ? _GEN_1666 : dirty_129; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1923 = ~_GEN_767 ? _GEN_1667 : dirty_130; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1924 = ~_GEN_767 ? _GEN_1668 : dirty_131; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1925 = ~_GEN_767 ? _GEN_1669 : dirty_132; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1926 = ~_GEN_767 ? _GEN_1670 : dirty_133; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1927 = ~_GEN_767 ? _GEN_1671 : dirty_134; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1928 = ~_GEN_767 ? _GEN_1672 : dirty_135; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1929 = ~_GEN_767 ? _GEN_1673 : dirty_136; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1930 = ~_GEN_767 ? _GEN_1674 : dirty_137; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1931 = ~_GEN_767 ? _GEN_1675 : dirty_138; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1932 = ~_GEN_767 ? _GEN_1676 : dirty_139; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1933 = ~_GEN_767 ? _GEN_1677 : dirty_140; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1934 = ~_GEN_767 ? _GEN_1678 : dirty_141; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1935 = ~_GEN_767 ? _GEN_1679 : dirty_142; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1936 = ~_GEN_767 ? _GEN_1680 : dirty_143; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1937 = ~_GEN_767 ? _GEN_1681 : dirty_144; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1938 = ~_GEN_767 ? _GEN_1682 : dirty_145; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1939 = ~_GEN_767 ? _GEN_1683 : dirty_146; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1940 = ~_GEN_767 ? _GEN_1684 : dirty_147; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1941 = ~_GEN_767 ? _GEN_1685 : dirty_148; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1942 = ~_GEN_767 ? _GEN_1686 : dirty_149; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1943 = ~_GEN_767 ? _GEN_1687 : dirty_150; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1944 = ~_GEN_767 ? _GEN_1688 : dirty_151; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1945 = ~_GEN_767 ? _GEN_1689 : dirty_152; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1946 = ~_GEN_767 ? _GEN_1690 : dirty_153; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1947 = ~_GEN_767 ? _GEN_1691 : dirty_154; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1948 = ~_GEN_767 ? _GEN_1692 : dirty_155; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1949 = ~_GEN_767 ? _GEN_1693 : dirty_156; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1950 = ~_GEN_767 ? _GEN_1694 : dirty_157; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1951 = ~_GEN_767 ? _GEN_1695 : dirty_158; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1952 = ~_GEN_767 ? _GEN_1696 : dirty_159; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1953 = ~_GEN_767 ? _GEN_1697 : dirty_160; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1954 = ~_GEN_767 ? _GEN_1698 : dirty_161; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1955 = ~_GEN_767 ? _GEN_1699 : dirty_162; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1956 = ~_GEN_767 ? _GEN_1700 : dirty_163; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1957 = ~_GEN_767 ? _GEN_1701 : dirty_164; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1958 = ~_GEN_767 ? _GEN_1702 : dirty_165; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1959 = ~_GEN_767 ? _GEN_1703 : dirty_166; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1960 = ~_GEN_767 ? _GEN_1704 : dirty_167; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1961 = ~_GEN_767 ? _GEN_1705 : dirty_168; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1962 = ~_GEN_767 ? _GEN_1706 : dirty_169; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1963 = ~_GEN_767 ? _GEN_1707 : dirty_170; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1964 = ~_GEN_767 ? _GEN_1708 : dirty_171; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1965 = ~_GEN_767 ? _GEN_1709 : dirty_172; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1966 = ~_GEN_767 ? _GEN_1710 : dirty_173; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1967 = ~_GEN_767 ? _GEN_1711 : dirty_174; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1968 = ~_GEN_767 ? _GEN_1712 : dirty_175; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1969 = ~_GEN_767 ? _GEN_1713 : dirty_176; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1970 = ~_GEN_767 ? _GEN_1714 : dirty_177; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1971 = ~_GEN_767 ? _GEN_1715 : dirty_178; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1972 = ~_GEN_767 ? _GEN_1716 : dirty_179; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1973 = ~_GEN_767 ? _GEN_1717 : dirty_180; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1974 = ~_GEN_767 ? _GEN_1718 : dirty_181; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1975 = ~_GEN_767 ? _GEN_1719 : dirty_182; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1976 = ~_GEN_767 ? _GEN_1720 : dirty_183; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1977 = ~_GEN_767 ? _GEN_1721 : dirty_184; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1978 = ~_GEN_767 ? _GEN_1722 : dirty_185; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1979 = ~_GEN_767 ? _GEN_1723 : dirty_186; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1980 = ~_GEN_767 ? _GEN_1724 : dirty_187; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1981 = ~_GEN_767 ? _GEN_1725 : dirty_188; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1982 = ~_GEN_767 ? _GEN_1726 : dirty_189; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1983 = ~_GEN_767 ? _GEN_1727 : dirty_190; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1984 = ~_GEN_767 ? _GEN_1728 : dirty_191; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1985 = ~_GEN_767 ? _GEN_1729 : dirty_192; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1986 = ~_GEN_767 ? _GEN_1730 : dirty_193; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1987 = ~_GEN_767 ? _GEN_1731 : dirty_194; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1988 = ~_GEN_767 ? _GEN_1732 : dirty_195; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1989 = ~_GEN_767 ? _GEN_1733 : dirty_196; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1990 = ~_GEN_767 ? _GEN_1734 : dirty_197; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1991 = ~_GEN_767 ? _GEN_1735 : dirty_198; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1992 = ~_GEN_767 ? _GEN_1736 : dirty_199; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1993 = ~_GEN_767 ? _GEN_1737 : dirty_200; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1994 = ~_GEN_767 ? _GEN_1738 : dirty_201; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1995 = ~_GEN_767 ? _GEN_1739 : dirty_202; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1996 = ~_GEN_767 ? _GEN_1740 : dirty_203; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1997 = ~_GEN_767 ? _GEN_1741 : dirty_204; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1998 = ~_GEN_767 ? _GEN_1742 : dirty_205; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_1999 = ~_GEN_767 ? _GEN_1743 : dirty_206; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2000 = ~_GEN_767 ? _GEN_1744 : dirty_207; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2001 = ~_GEN_767 ? _GEN_1745 : dirty_208; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2002 = ~_GEN_767 ? _GEN_1746 : dirty_209; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2003 = ~_GEN_767 ? _GEN_1747 : dirty_210; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2004 = ~_GEN_767 ? _GEN_1748 : dirty_211; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2005 = ~_GEN_767 ? _GEN_1749 : dirty_212; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2006 = ~_GEN_767 ? _GEN_1750 : dirty_213; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2007 = ~_GEN_767 ? _GEN_1751 : dirty_214; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2008 = ~_GEN_767 ? _GEN_1752 : dirty_215; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2009 = ~_GEN_767 ? _GEN_1753 : dirty_216; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2010 = ~_GEN_767 ? _GEN_1754 : dirty_217; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2011 = ~_GEN_767 ? _GEN_1755 : dirty_218; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2012 = ~_GEN_767 ? _GEN_1756 : dirty_219; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2013 = ~_GEN_767 ? _GEN_1757 : dirty_220; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2014 = ~_GEN_767 ? _GEN_1758 : dirty_221; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2015 = ~_GEN_767 ? _GEN_1759 : dirty_222; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2016 = ~_GEN_767 ? _GEN_1760 : dirty_223; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2017 = ~_GEN_767 ? _GEN_1761 : dirty_224; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2018 = ~_GEN_767 ? _GEN_1762 : dirty_225; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2019 = ~_GEN_767 ? _GEN_1763 : dirty_226; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2020 = ~_GEN_767 ? _GEN_1764 : dirty_227; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2021 = ~_GEN_767 ? _GEN_1765 : dirty_228; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2022 = ~_GEN_767 ? _GEN_1766 : dirty_229; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2023 = ~_GEN_767 ? _GEN_1767 : dirty_230; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2024 = ~_GEN_767 ? _GEN_1768 : dirty_231; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2025 = ~_GEN_767 ? _GEN_1769 : dirty_232; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2026 = ~_GEN_767 ? _GEN_1770 : dirty_233; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2027 = ~_GEN_767 ? _GEN_1771 : dirty_234; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2028 = ~_GEN_767 ? _GEN_1772 : dirty_235; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2029 = ~_GEN_767 ? _GEN_1773 : dirty_236; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2030 = ~_GEN_767 ? _GEN_1774 : dirty_237; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2031 = ~_GEN_767 ? _GEN_1775 : dirty_238; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2032 = ~_GEN_767 ? _GEN_1776 : dirty_239; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2033 = ~_GEN_767 ? _GEN_1777 : dirty_240; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2034 = ~_GEN_767 ? _GEN_1778 : dirty_241; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2035 = ~_GEN_767 ? _GEN_1779 : dirty_242; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2036 = ~_GEN_767 ? _GEN_1780 : dirty_243; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2037 = ~_GEN_767 ? _GEN_1781 : dirty_244; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2038 = ~_GEN_767 ? _GEN_1782 : dirty_245; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2039 = ~_GEN_767 ? _GEN_1783 : dirty_246; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2040 = ~_GEN_767 ? _GEN_1784 : dirty_247; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2041 = ~_GEN_767 ? _GEN_1785 : dirty_248; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2042 = ~_GEN_767 ? _GEN_1786 : dirty_249; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2043 = ~_GEN_767 ? _GEN_1787 : dirty_250; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2044 = ~_GEN_767 ? _GEN_1788 : dirty_251; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2045 = ~_GEN_767 ? _GEN_1789 : dirty_252; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2046 = ~_GEN_767 ? _GEN_1790 : dirty_253; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2047 = ~_GEN_767 ? _GEN_1791 : dirty_254; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire  _GEN_2048 = ~_GEN_767 ? _GEN_1792 : dirty_255; // @[Dcache.scala 139:34 Dcache.scala 18:24]
  wire [2:0] _GEN_2049 = cache_dirty ? 3'h2 : 3'h4; // @[Dcache.scala 144:31 Dcache.scala 145:15 Dcache.scala 148:15]
  wire  _GEN_2818 = cache_hit | data_ready; // @[Dcache.scala 131:24 Dcache.scala 135:27 Dcache.scala 46:28]
  wire  _T_3 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_3080 = 8'h1 == req_index ? offset_1 : offset_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3081 = 8'h2 == req_index ? offset_2 : _GEN_3080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3082 = 8'h3 == req_index ? offset_3 : _GEN_3081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3083 = 8'h4 == req_index ? offset_4 : _GEN_3082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3084 = 8'h5 == req_index ? offset_5 : _GEN_3083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3085 = 8'h6 == req_index ? offset_6 : _GEN_3084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3086 = 8'h7 == req_index ? offset_7 : _GEN_3085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3087 = 8'h8 == req_index ? offset_8 : _GEN_3086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3088 = 8'h9 == req_index ? offset_9 : _GEN_3087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3089 = 8'ha == req_index ? offset_10 : _GEN_3088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3090 = 8'hb == req_index ? offset_11 : _GEN_3089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3091 = 8'hc == req_index ? offset_12 : _GEN_3090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3092 = 8'hd == req_index ? offset_13 : _GEN_3091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3093 = 8'he == req_index ? offset_14 : _GEN_3092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3094 = 8'hf == req_index ? offset_15 : _GEN_3093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3095 = 8'h10 == req_index ? offset_16 : _GEN_3094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3096 = 8'h11 == req_index ? offset_17 : _GEN_3095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3097 = 8'h12 == req_index ? offset_18 : _GEN_3096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3098 = 8'h13 == req_index ? offset_19 : _GEN_3097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3099 = 8'h14 == req_index ? offset_20 : _GEN_3098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3100 = 8'h15 == req_index ? offset_21 : _GEN_3099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3101 = 8'h16 == req_index ? offset_22 : _GEN_3100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3102 = 8'h17 == req_index ? offset_23 : _GEN_3101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3103 = 8'h18 == req_index ? offset_24 : _GEN_3102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3104 = 8'h19 == req_index ? offset_25 : _GEN_3103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3105 = 8'h1a == req_index ? offset_26 : _GEN_3104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3106 = 8'h1b == req_index ? offset_27 : _GEN_3105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3107 = 8'h1c == req_index ? offset_28 : _GEN_3106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3108 = 8'h1d == req_index ? offset_29 : _GEN_3107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3109 = 8'h1e == req_index ? offset_30 : _GEN_3108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3110 = 8'h1f == req_index ? offset_31 : _GEN_3109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3111 = 8'h20 == req_index ? offset_32 : _GEN_3110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3112 = 8'h21 == req_index ? offset_33 : _GEN_3111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3113 = 8'h22 == req_index ? offset_34 : _GEN_3112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3114 = 8'h23 == req_index ? offset_35 : _GEN_3113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3115 = 8'h24 == req_index ? offset_36 : _GEN_3114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3116 = 8'h25 == req_index ? offset_37 : _GEN_3115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3117 = 8'h26 == req_index ? offset_38 : _GEN_3116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3118 = 8'h27 == req_index ? offset_39 : _GEN_3117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3119 = 8'h28 == req_index ? offset_40 : _GEN_3118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3120 = 8'h29 == req_index ? offset_41 : _GEN_3119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3121 = 8'h2a == req_index ? offset_42 : _GEN_3120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3122 = 8'h2b == req_index ? offset_43 : _GEN_3121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3123 = 8'h2c == req_index ? offset_44 : _GEN_3122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3124 = 8'h2d == req_index ? offset_45 : _GEN_3123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3125 = 8'h2e == req_index ? offset_46 : _GEN_3124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3126 = 8'h2f == req_index ? offset_47 : _GEN_3125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3127 = 8'h30 == req_index ? offset_48 : _GEN_3126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3128 = 8'h31 == req_index ? offset_49 : _GEN_3127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3129 = 8'h32 == req_index ? offset_50 : _GEN_3128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3130 = 8'h33 == req_index ? offset_51 : _GEN_3129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3131 = 8'h34 == req_index ? offset_52 : _GEN_3130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3132 = 8'h35 == req_index ? offset_53 : _GEN_3131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3133 = 8'h36 == req_index ? offset_54 : _GEN_3132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3134 = 8'h37 == req_index ? offset_55 : _GEN_3133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3135 = 8'h38 == req_index ? offset_56 : _GEN_3134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3136 = 8'h39 == req_index ? offset_57 : _GEN_3135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3137 = 8'h3a == req_index ? offset_58 : _GEN_3136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3138 = 8'h3b == req_index ? offset_59 : _GEN_3137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3139 = 8'h3c == req_index ? offset_60 : _GEN_3138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3140 = 8'h3d == req_index ? offset_61 : _GEN_3139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3141 = 8'h3e == req_index ? offset_62 : _GEN_3140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3142 = 8'h3f == req_index ? offset_63 : _GEN_3141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3143 = 8'h40 == req_index ? offset_64 : _GEN_3142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3144 = 8'h41 == req_index ? offset_65 : _GEN_3143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3145 = 8'h42 == req_index ? offset_66 : _GEN_3144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3146 = 8'h43 == req_index ? offset_67 : _GEN_3145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3147 = 8'h44 == req_index ? offset_68 : _GEN_3146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3148 = 8'h45 == req_index ? offset_69 : _GEN_3147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3149 = 8'h46 == req_index ? offset_70 : _GEN_3148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3150 = 8'h47 == req_index ? offset_71 : _GEN_3149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3151 = 8'h48 == req_index ? offset_72 : _GEN_3150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3152 = 8'h49 == req_index ? offset_73 : _GEN_3151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3153 = 8'h4a == req_index ? offset_74 : _GEN_3152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3154 = 8'h4b == req_index ? offset_75 : _GEN_3153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3155 = 8'h4c == req_index ? offset_76 : _GEN_3154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3156 = 8'h4d == req_index ? offset_77 : _GEN_3155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3157 = 8'h4e == req_index ? offset_78 : _GEN_3156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3158 = 8'h4f == req_index ? offset_79 : _GEN_3157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3159 = 8'h50 == req_index ? offset_80 : _GEN_3158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3160 = 8'h51 == req_index ? offset_81 : _GEN_3159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3161 = 8'h52 == req_index ? offset_82 : _GEN_3160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3162 = 8'h53 == req_index ? offset_83 : _GEN_3161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3163 = 8'h54 == req_index ? offset_84 : _GEN_3162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3164 = 8'h55 == req_index ? offset_85 : _GEN_3163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3165 = 8'h56 == req_index ? offset_86 : _GEN_3164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3166 = 8'h57 == req_index ? offset_87 : _GEN_3165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3167 = 8'h58 == req_index ? offset_88 : _GEN_3166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3168 = 8'h59 == req_index ? offset_89 : _GEN_3167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3169 = 8'h5a == req_index ? offset_90 : _GEN_3168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3170 = 8'h5b == req_index ? offset_91 : _GEN_3169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3171 = 8'h5c == req_index ? offset_92 : _GEN_3170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3172 = 8'h5d == req_index ? offset_93 : _GEN_3171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3173 = 8'h5e == req_index ? offset_94 : _GEN_3172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3174 = 8'h5f == req_index ? offset_95 : _GEN_3173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3175 = 8'h60 == req_index ? offset_96 : _GEN_3174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3176 = 8'h61 == req_index ? offset_97 : _GEN_3175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3177 = 8'h62 == req_index ? offset_98 : _GEN_3176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3178 = 8'h63 == req_index ? offset_99 : _GEN_3177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3179 = 8'h64 == req_index ? offset_100 : _GEN_3178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3180 = 8'h65 == req_index ? offset_101 : _GEN_3179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3181 = 8'h66 == req_index ? offset_102 : _GEN_3180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3182 = 8'h67 == req_index ? offset_103 : _GEN_3181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3183 = 8'h68 == req_index ? offset_104 : _GEN_3182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3184 = 8'h69 == req_index ? offset_105 : _GEN_3183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3185 = 8'h6a == req_index ? offset_106 : _GEN_3184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3186 = 8'h6b == req_index ? offset_107 : _GEN_3185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3187 = 8'h6c == req_index ? offset_108 : _GEN_3186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3188 = 8'h6d == req_index ? offset_109 : _GEN_3187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3189 = 8'h6e == req_index ? offset_110 : _GEN_3188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3190 = 8'h6f == req_index ? offset_111 : _GEN_3189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3191 = 8'h70 == req_index ? offset_112 : _GEN_3190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3192 = 8'h71 == req_index ? offset_113 : _GEN_3191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3193 = 8'h72 == req_index ? offset_114 : _GEN_3192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3194 = 8'h73 == req_index ? offset_115 : _GEN_3193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3195 = 8'h74 == req_index ? offset_116 : _GEN_3194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3196 = 8'h75 == req_index ? offset_117 : _GEN_3195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3197 = 8'h76 == req_index ? offset_118 : _GEN_3196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3198 = 8'h77 == req_index ? offset_119 : _GEN_3197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3199 = 8'h78 == req_index ? offset_120 : _GEN_3198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3200 = 8'h79 == req_index ? offset_121 : _GEN_3199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3201 = 8'h7a == req_index ? offset_122 : _GEN_3200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3202 = 8'h7b == req_index ? offset_123 : _GEN_3201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3203 = 8'h7c == req_index ? offset_124 : _GEN_3202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3204 = 8'h7d == req_index ? offset_125 : _GEN_3203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3205 = 8'h7e == req_index ? offset_126 : _GEN_3204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3206 = 8'h7f == req_index ? offset_127 : _GEN_3205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3207 = 8'h80 == req_index ? offset_128 : _GEN_3206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3208 = 8'h81 == req_index ? offset_129 : _GEN_3207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3209 = 8'h82 == req_index ? offset_130 : _GEN_3208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3210 = 8'h83 == req_index ? offset_131 : _GEN_3209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3211 = 8'h84 == req_index ? offset_132 : _GEN_3210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3212 = 8'h85 == req_index ? offset_133 : _GEN_3211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3213 = 8'h86 == req_index ? offset_134 : _GEN_3212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3214 = 8'h87 == req_index ? offset_135 : _GEN_3213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3215 = 8'h88 == req_index ? offset_136 : _GEN_3214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3216 = 8'h89 == req_index ? offset_137 : _GEN_3215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3217 = 8'h8a == req_index ? offset_138 : _GEN_3216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3218 = 8'h8b == req_index ? offset_139 : _GEN_3217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3219 = 8'h8c == req_index ? offset_140 : _GEN_3218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3220 = 8'h8d == req_index ? offset_141 : _GEN_3219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3221 = 8'h8e == req_index ? offset_142 : _GEN_3220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3222 = 8'h8f == req_index ? offset_143 : _GEN_3221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3223 = 8'h90 == req_index ? offset_144 : _GEN_3222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3224 = 8'h91 == req_index ? offset_145 : _GEN_3223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3225 = 8'h92 == req_index ? offset_146 : _GEN_3224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3226 = 8'h93 == req_index ? offset_147 : _GEN_3225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3227 = 8'h94 == req_index ? offset_148 : _GEN_3226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3228 = 8'h95 == req_index ? offset_149 : _GEN_3227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3229 = 8'h96 == req_index ? offset_150 : _GEN_3228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3230 = 8'h97 == req_index ? offset_151 : _GEN_3229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3231 = 8'h98 == req_index ? offset_152 : _GEN_3230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3232 = 8'h99 == req_index ? offset_153 : _GEN_3231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3233 = 8'h9a == req_index ? offset_154 : _GEN_3232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3234 = 8'h9b == req_index ? offset_155 : _GEN_3233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3235 = 8'h9c == req_index ? offset_156 : _GEN_3234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3236 = 8'h9d == req_index ? offset_157 : _GEN_3235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3237 = 8'h9e == req_index ? offset_158 : _GEN_3236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3238 = 8'h9f == req_index ? offset_159 : _GEN_3237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3239 = 8'ha0 == req_index ? offset_160 : _GEN_3238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3240 = 8'ha1 == req_index ? offset_161 : _GEN_3239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3241 = 8'ha2 == req_index ? offset_162 : _GEN_3240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3242 = 8'ha3 == req_index ? offset_163 : _GEN_3241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3243 = 8'ha4 == req_index ? offset_164 : _GEN_3242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3244 = 8'ha5 == req_index ? offset_165 : _GEN_3243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3245 = 8'ha6 == req_index ? offset_166 : _GEN_3244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3246 = 8'ha7 == req_index ? offset_167 : _GEN_3245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3247 = 8'ha8 == req_index ? offset_168 : _GEN_3246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3248 = 8'ha9 == req_index ? offset_169 : _GEN_3247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3249 = 8'haa == req_index ? offset_170 : _GEN_3248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3250 = 8'hab == req_index ? offset_171 : _GEN_3249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3251 = 8'hac == req_index ? offset_172 : _GEN_3250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3252 = 8'had == req_index ? offset_173 : _GEN_3251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3253 = 8'hae == req_index ? offset_174 : _GEN_3252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3254 = 8'haf == req_index ? offset_175 : _GEN_3253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3255 = 8'hb0 == req_index ? offset_176 : _GEN_3254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3256 = 8'hb1 == req_index ? offset_177 : _GEN_3255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3257 = 8'hb2 == req_index ? offset_178 : _GEN_3256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3258 = 8'hb3 == req_index ? offset_179 : _GEN_3257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3259 = 8'hb4 == req_index ? offset_180 : _GEN_3258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3260 = 8'hb5 == req_index ? offset_181 : _GEN_3259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3261 = 8'hb6 == req_index ? offset_182 : _GEN_3260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3262 = 8'hb7 == req_index ? offset_183 : _GEN_3261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3263 = 8'hb8 == req_index ? offset_184 : _GEN_3262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3264 = 8'hb9 == req_index ? offset_185 : _GEN_3263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3265 = 8'hba == req_index ? offset_186 : _GEN_3264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3266 = 8'hbb == req_index ? offset_187 : _GEN_3265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3267 = 8'hbc == req_index ? offset_188 : _GEN_3266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3268 = 8'hbd == req_index ? offset_189 : _GEN_3267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3269 = 8'hbe == req_index ? offset_190 : _GEN_3268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3270 = 8'hbf == req_index ? offset_191 : _GEN_3269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3271 = 8'hc0 == req_index ? offset_192 : _GEN_3270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3272 = 8'hc1 == req_index ? offset_193 : _GEN_3271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3273 = 8'hc2 == req_index ? offset_194 : _GEN_3272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3274 = 8'hc3 == req_index ? offset_195 : _GEN_3273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3275 = 8'hc4 == req_index ? offset_196 : _GEN_3274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3276 = 8'hc5 == req_index ? offset_197 : _GEN_3275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3277 = 8'hc6 == req_index ? offset_198 : _GEN_3276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3278 = 8'hc7 == req_index ? offset_199 : _GEN_3277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3279 = 8'hc8 == req_index ? offset_200 : _GEN_3278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3280 = 8'hc9 == req_index ? offset_201 : _GEN_3279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3281 = 8'hca == req_index ? offset_202 : _GEN_3280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3282 = 8'hcb == req_index ? offset_203 : _GEN_3281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3283 = 8'hcc == req_index ? offset_204 : _GEN_3282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3284 = 8'hcd == req_index ? offset_205 : _GEN_3283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3285 = 8'hce == req_index ? offset_206 : _GEN_3284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3286 = 8'hcf == req_index ? offset_207 : _GEN_3285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3287 = 8'hd0 == req_index ? offset_208 : _GEN_3286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3288 = 8'hd1 == req_index ? offset_209 : _GEN_3287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3289 = 8'hd2 == req_index ? offset_210 : _GEN_3288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3290 = 8'hd3 == req_index ? offset_211 : _GEN_3289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3291 = 8'hd4 == req_index ? offset_212 : _GEN_3290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3292 = 8'hd5 == req_index ? offset_213 : _GEN_3291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3293 = 8'hd6 == req_index ? offset_214 : _GEN_3292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3294 = 8'hd7 == req_index ? offset_215 : _GEN_3293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3295 = 8'hd8 == req_index ? offset_216 : _GEN_3294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3296 = 8'hd9 == req_index ? offset_217 : _GEN_3295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3297 = 8'hda == req_index ? offset_218 : _GEN_3296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3298 = 8'hdb == req_index ? offset_219 : _GEN_3297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3299 = 8'hdc == req_index ? offset_220 : _GEN_3298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3300 = 8'hdd == req_index ? offset_221 : _GEN_3299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3301 = 8'hde == req_index ? offset_222 : _GEN_3300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3302 = 8'hdf == req_index ? offset_223 : _GEN_3301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3303 = 8'he0 == req_index ? offset_224 : _GEN_3302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3304 = 8'he1 == req_index ? offset_225 : _GEN_3303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3305 = 8'he2 == req_index ? offset_226 : _GEN_3304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3306 = 8'he3 == req_index ? offset_227 : _GEN_3305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3307 = 8'he4 == req_index ? offset_228 : _GEN_3306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3308 = 8'he5 == req_index ? offset_229 : _GEN_3307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3309 = 8'he6 == req_index ? offset_230 : _GEN_3308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3310 = 8'he7 == req_index ? offset_231 : _GEN_3309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3311 = 8'he8 == req_index ? offset_232 : _GEN_3310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3312 = 8'he9 == req_index ? offset_233 : _GEN_3311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3313 = 8'hea == req_index ? offset_234 : _GEN_3312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3314 = 8'heb == req_index ? offset_235 : _GEN_3313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3315 = 8'hec == req_index ? offset_236 : _GEN_3314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3316 = 8'hed == req_index ? offset_237 : _GEN_3315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3317 = 8'hee == req_index ? offset_238 : _GEN_3316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3318 = 8'hef == req_index ? offset_239 : _GEN_3317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3319 = 8'hf0 == req_index ? offset_240 : _GEN_3318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3320 = 8'hf1 == req_index ? offset_241 : _GEN_3319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3321 = 8'hf2 == req_index ? offset_242 : _GEN_3320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3322 = 8'hf3 == req_index ? offset_243 : _GEN_3321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3323 = 8'hf4 == req_index ? offset_244 : _GEN_3322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3324 = 8'hf5 == req_index ? offset_245 : _GEN_3323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3325 = 8'hf6 == req_index ? offset_246 : _GEN_3324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3326 = 8'hf7 == req_index ? offset_247 : _GEN_3325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3327 = 8'hf8 == req_index ? offset_248 : _GEN_3326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3328 = 8'hf9 == req_index ? offset_249 : _GEN_3327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3329 = 8'hfa == req_index ? offset_250 : _GEN_3328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3330 = 8'hfb == req_index ? offset_251 : _GEN_3329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3331 = 8'hfc == req_index ? offset_252 : _GEN_3330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3332 = 8'hfd == req_index ? offset_253 : _GEN_3331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3333 = 8'hfe == req_index ? offset_254 : _GEN_3332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3334 = 8'hff == req_index ? offset_255 : _GEN_3333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _data_addr_T = {_GEN_255,req_index,_GEN_3334}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_3335 = io_out_data_ready ? 3'h3 : 3'h2; // @[Dcache.scala 159:31 Dcache.scala 160:25 Dcache.scala 165:19]
  wire  _GEN_3336 = io_out_data_ready ? 1'h0 : 1'h1; // @[Dcache.scala 159:31 Dcache.scala 161:25 Dcache.scala 157:21]
  wire  _T_4 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_6 = ~cache_fill; // @[Dcache.scala 174:13]
  wire [2:0] _GEN_3337 = ~cache_fill ? 3'h4 : 3'h5; // @[Dcache.scala 174:26 Dcache.scala 175:21 Dcache.scala 184:15]
  wire [31:0] _GEN_3338 = ~cache_fill ? io_dmem_data_addr : 32'h0; // @[Dcache.scala 174:26 Dcache.scala 176:21]
  wire [127:0] _cache_wdata_T_5 = {valid_wdata,io_out_data_read[63:0]}; // @[Cat.scala 30:58]
  wire [127:0] _cache_wdata_T_6 = {io_out_data_read[127:64],valid_wdata}; // @[Cat.scala 30:58]
  wire [127:0] _cache_wdata_T_7 = req_offset[3] ? _cache_wdata_T_5 : _cache_wdata_T_6; // @[Dcache.scala 189:44]
  wire [127:0] _cache_wdata_T_8 = io_dmem_data_req ? _cache_wdata_T_7 : io_out_data_read; // @[Dcache.scala 189:27]
  wire  _GEN_3344 = io_out_data_ready | cache_fill; // @[Dcache.scala 186:29 Dcache.scala 187:21 Dcache.scala 116:28]
  wire  _GEN_3345 = io_out_data_ready | cache_wen; // @[Dcache.scala 186:29 Dcache.scala 188:21 Dcache.scala 117:28]
  wire [127:0] _GEN_3346 = io_out_data_ready ? _cache_wdata_T_8 : cache_wdata; // @[Dcache.scala 186:29 Dcache.scala 189:21 Dcache.scala 118:28]
  wire [127:0] _GEN_3347 = io_out_data_ready ? 128'hffffffffffffffffffffffffffffffff : cache_strb; // @[Dcache.scala 186:29 Dcache.scala 190:21 Dcache.scala 119:28]
  wire  _GEN_3348 = io_out_data_ready ? 1'h0 : _T_6; // @[Dcache.scala 186:29 Dcache.scala 191:21]
  wire  _T_7 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_4373 = _T_7 ? 1'h0 : cache_fill; // @[Conditional.scala 39:67 Dcache.scala 196:25 Dcache.scala 116:28]
  wire  _GEN_4374 = _T_7 | data_ready; // @[Conditional.scala 39:67 Dcache.scala 197:25 Dcache.scala 46:28]
  wire  _GEN_4375 = _T_7 ? 1'h0 : cache_wen; // @[Conditional.scala 39:67 Dcache.scala 198:25 Dcache.scala 117:28]
  wire  _GEN_4376 = _T_7 ? _GEN_769 : valid_0; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4377 = _T_7 ? _GEN_770 : valid_1; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4378 = _T_7 ? _GEN_771 : valid_2; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4379 = _T_7 ? _GEN_772 : valid_3; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4380 = _T_7 ? _GEN_773 : valid_4; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4381 = _T_7 ? _GEN_774 : valid_5; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4382 = _T_7 ? _GEN_775 : valid_6; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4383 = _T_7 ? _GEN_776 : valid_7; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4384 = _T_7 ? _GEN_777 : valid_8; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4385 = _T_7 ? _GEN_778 : valid_9; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4386 = _T_7 ? _GEN_779 : valid_10; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4387 = _T_7 ? _GEN_780 : valid_11; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4388 = _T_7 ? _GEN_781 : valid_12; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4389 = _T_7 ? _GEN_782 : valid_13; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4390 = _T_7 ? _GEN_783 : valid_14; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4391 = _T_7 ? _GEN_784 : valid_15; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4392 = _T_7 ? _GEN_785 : valid_16; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4393 = _T_7 ? _GEN_786 : valid_17; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4394 = _T_7 ? _GEN_787 : valid_18; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4395 = _T_7 ? _GEN_788 : valid_19; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4396 = _T_7 ? _GEN_789 : valid_20; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4397 = _T_7 ? _GEN_790 : valid_21; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4398 = _T_7 ? _GEN_791 : valid_22; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4399 = _T_7 ? _GEN_792 : valid_23; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4400 = _T_7 ? _GEN_793 : valid_24; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4401 = _T_7 ? _GEN_794 : valid_25; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4402 = _T_7 ? _GEN_795 : valid_26; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4403 = _T_7 ? _GEN_796 : valid_27; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4404 = _T_7 ? _GEN_797 : valid_28; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4405 = _T_7 ? _GEN_798 : valid_29; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4406 = _T_7 ? _GEN_799 : valid_30; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4407 = _T_7 ? _GEN_800 : valid_31; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4408 = _T_7 ? _GEN_801 : valid_32; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4409 = _T_7 ? _GEN_802 : valid_33; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4410 = _T_7 ? _GEN_803 : valid_34; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4411 = _T_7 ? _GEN_804 : valid_35; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4412 = _T_7 ? _GEN_805 : valid_36; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4413 = _T_7 ? _GEN_806 : valid_37; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4414 = _T_7 ? _GEN_807 : valid_38; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4415 = _T_7 ? _GEN_808 : valid_39; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4416 = _T_7 ? _GEN_809 : valid_40; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4417 = _T_7 ? _GEN_810 : valid_41; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4418 = _T_7 ? _GEN_811 : valid_42; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4419 = _T_7 ? _GEN_812 : valid_43; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4420 = _T_7 ? _GEN_813 : valid_44; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4421 = _T_7 ? _GEN_814 : valid_45; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4422 = _T_7 ? _GEN_815 : valid_46; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4423 = _T_7 ? _GEN_816 : valid_47; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4424 = _T_7 ? _GEN_817 : valid_48; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4425 = _T_7 ? _GEN_818 : valid_49; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4426 = _T_7 ? _GEN_819 : valid_50; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4427 = _T_7 ? _GEN_820 : valid_51; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4428 = _T_7 ? _GEN_821 : valid_52; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4429 = _T_7 ? _GEN_822 : valid_53; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4430 = _T_7 ? _GEN_823 : valid_54; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4431 = _T_7 ? _GEN_824 : valid_55; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4432 = _T_7 ? _GEN_825 : valid_56; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4433 = _T_7 ? _GEN_826 : valid_57; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4434 = _T_7 ? _GEN_827 : valid_58; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4435 = _T_7 ? _GEN_828 : valid_59; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4436 = _T_7 ? _GEN_829 : valid_60; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4437 = _T_7 ? _GEN_830 : valid_61; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4438 = _T_7 ? _GEN_831 : valid_62; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4439 = _T_7 ? _GEN_832 : valid_63; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4440 = _T_7 ? _GEN_833 : valid_64; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4441 = _T_7 ? _GEN_834 : valid_65; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4442 = _T_7 ? _GEN_835 : valid_66; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4443 = _T_7 ? _GEN_836 : valid_67; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4444 = _T_7 ? _GEN_837 : valid_68; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4445 = _T_7 ? _GEN_838 : valid_69; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4446 = _T_7 ? _GEN_839 : valid_70; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4447 = _T_7 ? _GEN_840 : valid_71; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4448 = _T_7 ? _GEN_841 : valid_72; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4449 = _T_7 ? _GEN_842 : valid_73; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4450 = _T_7 ? _GEN_843 : valid_74; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4451 = _T_7 ? _GEN_844 : valid_75; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4452 = _T_7 ? _GEN_845 : valid_76; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4453 = _T_7 ? _GEN_846 : valid_77; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4454 = _T_7 ? _GEN_847 : valid_78; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4455 = _T_7 ? _GEN_848 : valid_79; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4456 = _T_7 ? _GEN_849 : valid_80; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4457 = _T_7 ? _GEN_850 : valid_81; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4458 = _T_7 ? _GEN_851 : valid_82; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4459 = _T_7 ? _GEN_852 : valid_83; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4460 = _T_7 ? _GEN_853 : valid_84; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4461 = _T_7 ? _GEN_854 : valid_85; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4462 = _T_7 ? _GEN_855 : valid_86; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4463 = _T_7 ? _GEN_856 : valid_87; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4464 = _T_7 ? _GEN_857 : valid_88; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4465 = _T_7 ? _GEN_858 : valid_89; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4466 = _T_7 ? _GEN_859 : valid_90; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4467 = _T_7 ? _GEN_860 : valid_91; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4468 = _T_7 ? _GEN_861 : valid_92; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4469 = _T_7 ? _GEN_862 : valid_93; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4470 = _T_7 ? _GEN_863 : valid_94; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4471 = _T_7 ? _GEN_864 : valid_95; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4472 = _T_7 ? _GEN_865 : valid_96; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4473 = _T_7 ? _GEN_866 : valid_97; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4474 = _T_7 ? _GEN_867 : valid_98; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4475 = _T_7 ? _GEN_868 : valid_99; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4476 = _T_7 ? _GEN_869 : valid_100; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4477 = _T_7 ? _GEN_870 : valid_101; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4478 = _T_7 ? _GEN_871 : valid_102; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4479 = _T_7 ? _GEN_872 : valid_103; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4480 = _T_7 ? _GEN_873 : valid_104; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4481 = _T_7 ? _GEN_874 : valid_105; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4482 = _T_7 ? _GEN_875 : valid_106; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4483 = _T_7 ? _GEN_876 : valid_107; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4484 = _T_7 ? _GEN_877 : valid_108; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4485 = _T_7 ? _GEN_878 : valid_109; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4486 = _T_7 ? _GEN_879 : valid_110; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4487 = _T_7 ? _GEN_880 : valid_111; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4488 = _T_7 ? _GEN_881 : valid_112; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4489 = _T_7 ? _GEN_882 : valid_113; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4490 = _T_7 ? _GEN_883 : valid_114; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4491 = _T_7 ? _GEN_884 : valid_115; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4492 = _T_7 ? _GEN_885 : valid_116; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4493 = _T_7 ? _GEN_886 : valid_117; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4494 = _T_7 ? _GEN_887 : valid_118; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4495 = _T_7 ? _GEN_888 : valid_119; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4496 = _T_7 ? _GEN_889 : valid_120; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4497 = _T_7 ? _GEN_890 : valid_121; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4498 = _T_7 ? _GEN_891 : valid_122; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4499 = _T_7 ? _GEN_892 : valid_123; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4500 = _T_7 ? _GEN_893 : valid_124; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4501 = _T_7 ? _GEN_894 : valid_125; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4502 = _T_7 ? _GEN_895 : valid_126; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4503 = _T_7 ? _GEN_896 : valid_127; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4504 = _T_7 ? _GEN_897 : valid_128; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4505 = _T_7 ? _GEN_898 : valid_129; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4506 = _T_7 ? _GEN_899 : valid_130; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4507 = _T_7 ? _GEN_900 : valid_131; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4508 = _T_7 ? _GEN_901 : valid_132; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4509 = _T_7 ? _GEN_902 : valid_133; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4510 = _T_7 ? _GEN_903 : valid_134; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4511 = _T_7 ? _GEN_904 : valid_135; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4512 = _T_7 ? _GEN_905 : valid_136; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4513 = _T_7 ? _GEN_906 : valid_137; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4514 = _T_7 ? _GEN_907 : valid_138; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4515 = _T_7 ? _GEN_908 : valid_139; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4516 = _T_7 ? _GEN_909 : valid_140; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4517 = _T_7 ? _GEN_910 : valid_141; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4518 = _T_7 ? _GEN_911 : valid_142; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4519 = _T_7 ? _GEN_912 : valid_143; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4520 = _T_7 ? _GEN_913 : valid_144; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4521 = _T_7 ? _GEN_914 : valid_145; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4522 = _T_7 ? _GEN_915 : valid_146; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4523 = _T_7 ? _GEN_916 : valid_147; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4524 = _T_7 ? _GEN_917 : valid_148; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4525 = _T_7 ? _GEN_918 : valid_149; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4526 = _T_7 ? _GEN_919 : valid_150; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4527 = _T_7 ? _GEN_920 : valid_151; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4528 = _T_7 ? _GEN_921 : valid_152; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4529 = _T_7 ? _GEN_922 : valid_153; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4530 = _T_7 ? _GEN_923 : valid_154; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4531 = _T_7 ? _GEN_924 : valid_155; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4532 = _T_7 ? _GEN_925 : valid_156; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4533 = _T_7 ? _GEN_926 : valid_157; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4534 = _T_7 ? _GEN_927 : valid_158; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4535 = _T_7 ? _GEN_928 : valid_159; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4536 = _T_7 ? _GEN_929 : valid_160; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4537 = _T_7 ? _GEN_930 : valid_161; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4538 = _T_7 ? _GEN_931 : valid_162; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4539 = _T_7 ? _GEN_932 : valid_163; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4540 = _T_7 ? _GEN_933 : valid_164; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4541 = _T_7 ? _GEN_934 : valid_165; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4542 = _T_7 ? _GEN_935 : valid_166; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4543 = _T_7 ? _GEN_936 : valid_167; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4544 = _T_7 ? _GEN_937 : valid_168; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4545 = _T_7 ? _GEN_938 : valid_169; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4546 = _T_7 ? _GEN_939 : valid_170; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4547 = _T_7 ? _GEN_940 : valid_171; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4548 = _T_7 ? _GEN_941 : valid_172; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4549 = _T_7 ? _GEN_942 : valid_173; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4550 = _T_7 ? _GEN_943 : valid_174; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4551 = _T_7 ? _GEN_944 : valid_175; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4552 = _T_7 ? _GEN_945 : valid_176; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4553 = _T_7 ? _GEN_946 : valid_177; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4554 = _T_7 ? _GEN_947 : valid_178; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4555 = _T_7 ? _GEN_948 : valid_179; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4556 = _T_7 ? _GEN_949 : valid_180; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4557 = _T_7 ? _GEN_950 : valid_181; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4558 = _T_7 ? _GEN_951 : valid_182; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4559 = _T_7 ? _GEN_952 : valid_183; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4560 = _T_7 ? _GEN_953 : valid_184; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4561 = _T_7 ? _GEN_954 : valid_185; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4562 = _T_7 ? _GEN_955 : valid_186; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4563 = _T_7 ? _GEN_956 : valid_187; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4564 = _T_7 ? _GEN_957 : valid_188; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4565 = _T_7 ? _GEN_958 : valid_189; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4566 = _T_7 ? _GEN_959 : valid_190; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4567 = _T_7 ? _GEN_960 : valid_191; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4568 = _T_7 ? _GEN_961 : valid_192; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4569 = _T_7 ? _GEN_962 : valid_193; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4570 = _T_7 ? _GEN_963 : valid_194; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4571 = _T_7 ? _GEN_964 : valid_195; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4572 = _T_7 ? _GEN_965 : valid_196; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4573 = _T_7 ? _GEN_966 : valid_197; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4574 = _T_7 ? _GEN_967 : valid_198; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4575 = _T_7 ? _GEN_968 : valid_199; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4576 = _T_7 ? _GEN_969 : valid_200; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4577 = _T_7 ? _GEN_970 : valid_201; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4578 = _T_7 ? _GEN_971 : valid_202; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4579 = _T_7 ? _GEN_972 : valid_203; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4580 = _T_7 ? _GEN_973 : valid_204; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4581 = _T_7 ? _GEN_974 : valid_205; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4582 = _T_7 ? _GEN_975 : valid_206; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4583 = _T_7 ? _GEN_976 : valid_207; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4584 = _T_7 ? _GEN_977 : valid_208; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4585 = _T_7 ? _GEN_978 : valid_209; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4586 = _T_7 ? _GEN_979 : valid_210; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4587 = _T_7 ? _GEN_980 : valid_211; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4588 = _T_7 ? _GEN_981 : valid_212; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4589 = _T_7 ? _GEN_982 : valid_213; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4590 = _T_7 ? _GEN_983 : valid_214; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4591 = _T_7 ? _GEN_984 : valid_215; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4592 = _T_7 ? _GEN_985 : valid_216; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4593 = _T_7 ? _GEN_986 : valid_217; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4594 = _T_7 ? _GEN_987 : valid_218; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4595 = _T_7 ? _GEN_988 : valid_219; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4596 = _T_7 ? _GEN_989 : valid_220; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4597 = _T_7 ? _GEN_990 : valid_221; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4598 = _T_7 ? _GEN_991 : valid_222; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4599 = _T_7 ? _GEN_992 : valid_223; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4600 = _T_7 ? _GEN_993 : valid_224; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4601 = _T_7 ? _GEN_994 : valid_225; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4602 = _T_7 ? _GEN_995 : valid_226; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4603 = _T_7 ? _GEN_996 : valid_227; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4604 = _T_7 ? _GEN_997 : valid_228; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4605 = _T_7 ? _GEN_998 : valid_229; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4606 = _T_7 ? _GEN_999 : valid_230; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4607 = _T_7 ? _GEN_1000 : valid_231; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4608 = _T_7 ? _GEN_1001 : valid_232; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4609 = _T_7 ? _GEN_1002 : valid_233; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4610 = _T_7 ? _GEN_1003 : valid_234; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4611 = _T_7 ? _GEN_1004 : valid_235; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4612 = _T_7 ? _GEN_1005 : valid_236; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4613 = _T_7 ? _GEN_1006 : valid_237; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4614 = _T_7 ? _GEN_1007 : valid_238; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4615 = _T_7 ? _GEN_1008 : valid_239; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4616 = _T_7 ? _GEN_1009 : valid_240; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4617 = _T_7 ? _GEN_1010 : valid_241; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4618 = _T_7 ? _GEN_1011 : valid_242; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4619 = _T_7 ? _GEN_1012 : valid_243; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4620 = _T_7 ? _GEN_1013 : valid_244; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4621 = _T_7 ? _GEN_1014 : valid_245; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4622 = _T_7 ? _GEN_1015 : valid_246; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4623 = _T_7 ? _GEN_1016 : valid_247; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4624 = _T_7 ? _GEN_1017 : valid_248; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4625 = _T_7 ? _GEN_1018 : valid_249; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4626 = _T_7 ? _GEN_1019 : valid_250; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4627 = _T_7 ? _GEN_1020 : valid_251; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4628 = _T_7 ? _GEN_1021 : valid_252; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4629 = _T_7 ? _GEN_1022 : valid_253; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4630 = _T_7 ? _GEN_1023 : valid_254; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_4631 = _T_7 ? _GEN_1024 : valid_255; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire [19:0] _GEN_4632 = _T_7 ? _GEN_1025 : tag_0; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4633 = _T_7 ? _GEN_1026 : tag_1; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4634 = _T_7 ? _GEN_1027 : tag_2; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4635 = _T_7 ? _GEN_1028 : tag_3; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4636 = _T_7 ? _GEN_1029 : tag_4; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4637 = _T_7 ? _GEN_1030 : tag_5; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4638 = _T_7 ? _GEN_1031 : tag_6; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4639 = _T_7 ? _GEN_1032 : tag_7; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4640 = _T_7 ? _GEN_1033 : tag_8; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4641 = _T_7 ? _GEN_1034 : tag_9; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4642 = _T_7 ? _GEN_1035 : tag_10; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4643 = _T_7 ? _GEN_1036 : tag_11; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4644 = _T_7 ? _GEN_1037 : tag_12; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4645 = _T_7 ? _GEN_1038 : tag_13; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4646 = _T_7 ? _GEN_1039 : tag_14; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4647 = _T_7 ? _GEN_1040 : tag_15; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4648 = _T_7 ? _GEN_1041 : tag_16; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4649 = _T_7 ? _GEN_1042 : tag_17; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4650 = _T_7 ? _GEN_1043 : tag_18; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4651 = _T_7 ? _GEN_1044 : tag_19; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4652 = _T_7 ? _GEN_1045 : tag_20; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4653 = _T_7 ? _GEN_1046 : tag_21; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4654 = _T_7 ? _GEN_1047 : tag_22; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4655 = _T_7 ? _GEN_1048 : tag_23; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4656 = _T_7 ? _GEN_1049 : tag_24; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4657 = _T_7 ? _GEN_1050 : tag_25; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4658 = _T_7 ? _GEN_1051 : tag_26; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4659 = _T_7 ? _GEN_1052 : tag_27; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4660 = _T_7 ? _GEN_1053 : tag_28; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4661 = _T_7 ? _GEN_1054 : tag_29; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4662 = _T_7 ? _GEN_1055 : tag_30; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4663 = _T_7 ? _GEN_1056 : tag_31; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4664 = _T_7 ? _GEN_1057 : tag_32; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4665 = _T_7 ? _GEN_1058 : tag_33; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4666 = _T_7 ? _GEN_1059 : tag_34; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4667 = _T_7 ? _GEN_1060 : tag_35; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4668 = _T_7 ? _GEN_1061 : tag_36; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4669 = _T_7 ? _GEN_1062 : tag_37; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4670 = _T_7 ? _GEN_1063 : tag_38; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4671 = _T_7 ? _GEN_1064 : tag_39; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4672 = _T_7 ? _GEN_1065 : tag_40; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4673 = _T_7 ? _GEN_1066 : tag_41; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4674 = _T_7 ? _GEN_1067 : tag_42; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4675 = _T_7 ? _GEN_1068 : tag_43; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4676 = _T_7 ? _GEN_1069 : tag_44; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4677 = _T_7 ? _GEN_1070 : tag_45; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4678 = _T_7 ? _GEN_1071 : tag_46; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4679 = _T_7 ? _GEN_1072 : tag_47; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4680 = _T_7 ? _GEN_1073 : tag_48; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4681 = _T_7 ? _GEN_1074 : tag_49; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4682 = _T_7 ? _GEN_1075 : tag_50; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4683 = _T_7 ? _GEN_1076 : tag_51; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4684 = _T_7 ? _GEN_1077 : tag_52; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4685 = _T_7 ? _GEN_1078 : tag_53; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4686 = _T_7 ? _GEN_1079 : tag_54; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4687 = _T_7 ? _GEN_1080 : tag_55; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4688 = _T_7 ? _GEN_1081 : tag_56; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4689 = _T_7 ? _GEN_1082 : tag_57; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4690 = _T_7 ? _GEN_1083 : tag_58; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4691 = _T_7 ? _GEN_1084 : tag_59; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4692 = _T_7 ? _GEN_1085 : tag_60; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4693 = _T_7 ? _GEN_1086 : tag_61; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4694 = _T_7 ? _GEN_1087 : tag_62; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4695 = _T_7 ? _GEN_1088 : tag_63; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4696 = _T_7 ? _GEN_1089 : tag_64; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4697 = _T_7 ? _GEN_1090 : tag_65; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4698 = _T_7 ? _GEN_1091 : tag_66; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4699 = _T_7 ? _GEN_1092 : tag_67; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4700 = _T_7 ? _GEN_1093 : tag_68; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4701 = _T_7 ? _GEN_1094 : tag_69; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4702 = _T_7 ? _GEN_1095 : tag_70; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4703 = _T_7 ? _GEN_1096 : tag_71; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4704 = _T_7 ? _GEN_1097 : tag_72; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4705 = _T_7 ? _GEN_1098 : tag_73; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4706 = _T_7 ? _GEN_1099 : tag_74; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4707 = _T_7 ? _GEN_1100 : tag_75; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4708 = _T_7 ? _GEN_1101 : tag_76; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4709 = _T_7 ? _GEN_1102 : tag_77; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4710 = _T_7 ? _GEN_1103 : tag_78; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4711 = _T_7 ? _GEN_1104 : tag_79; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4712 = _T_7 ? _GEN_1105 : tag_80; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4713 = _T_7 ? _GEN_1106 : tag_81; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4714 = _T_7 ? _GEN_1107 : tag_82; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4715 = _T_7 ? _GEN_1108 : tag_83; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4716 = _T_7 ? _GEN_1109 : tag_84; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4717 = _T_7 ? _GEN_1110 : tag_85; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4718 = _T_7 ? _GEN_1111 : tag_86; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4719 = _T_7 ? _GEN_1112 : tag_87; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4720 = _T_7 ? _GEN_1113 : tag_88; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4721 = _T_7 ? _GEN_1114 : tag_89; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4722 = _T_7 ? _GEN_1115 : tag_90; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4723 = _T_7 ? _GEN_1116 : tag_91; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4724 = _T_7 ? _GEN_1117 : tag_92; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4725 = _T_7 ? _GEN_1118 : tag_93; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4726 = _T_7 ? _GEN_1119 : tag_94; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4727 = _T_7 ? _GEN_1120 : tag_95; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4728 = _T_7 ? _GEN_1121 : tag_96; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4729 = _T_7 ? _GEN_1122 : tag_97; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4730 = _T_7 ? _GEN_1123 : tag_98; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4731 = _T_7 ? _GEN_1124 : tag_99; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4732 = _T_7 ? _GEN_1125 : tag_100; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4733 = _T_7 ? _GEN_1126 : tag_101; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4734 = _T_7 ? _GEN_1127 : tag_102; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4735 = _T_7 ? _GEN_1128 : tag_103; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4736 = _T_7 ? _GEN_1129 : tag_104; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4737 = _T_7 ? _GEN_1130 : tag_105; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4738 = _T_7 ? _GEN_1131 : tag_106; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4739 = _T_7 ? _GEN_1132 : tag_107; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4740 = _T_7 ? _GEN_1133 : tag_108; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4741 = _T_7 ? _GEN_1134 : tag_109; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4742 = _T_7 ? _GEN_1135 : tag_110; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4743 = _T_7 ? _GEN_1136 : tag_111; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4744 = _T_7 ? _GEN_1137 : tag_112; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4745 = _T_7 ? _GEN_1138 : tag_113; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4746 = _T_7 ? _GEN_1139 : tag_114; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4747 = _T_7 ? _GEN_1140 : tag_115; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4748 = _T_7 ? _GEN_1141 : tag_116; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4749 = _T_7 ? _GEN_1142 : tag_117; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4750 = _T_7 ? _GEN_1143 : tag_118; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4751 = _T_7 ? _GEN_1144 : tag_119; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4752 = _T_7 ? _GEN_1145 : tag_120; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4753 = _T_7 ? _GEN_1146 : tag_121; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4754 = _T_7 ? _GEN_1147 : tag_122; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4755 = _T_7 ? _GEN_1148 : tag_123; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4756 = _T_7 ? _GEN_1149 : tag_124; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4757 = _T_7 ? _GEN_1150 : tag_125; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4758 = _T_7 ? _GEN_1151 : tag_126; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4759 = _T_7 ? _GEN_1152 : tag_127; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4760 = _T_7 ? _GEN_1153 : tag_128; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4761 = _T_7 ? _GEN_1154 : tag_129; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4762 = _T_7 ? _GEN_1155 : tag_130; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4763 = _T_7 ? _GEN_1156 : tag_131; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4764 = _T_7 ? _GEN_1157 : tag_132; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4765 = _T_7 ? _GEN_1158 : tag_133; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4766 = _T_7 ? _GEN_1159 : tag_134; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4767 = _T_7 ? _GEN_1160 : tag_135; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4768 = _T_7 ? _GEN_1161 : tag_136; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4769 = _T_7 ? _GEN_1162 : tag_137; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4770 = _T_7 ? _GEN_1163 : tag_138; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4771 = _T_7 ? _GEN_1164 : tag_139; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4772 = _T_7 ? _GEN_1165 : tag_140; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4773 = _T_7 ? _GEN_1166 : tag_141; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4774 = _T_7 ? _GEN_1167 : tag_142; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4775 = _T_7 ? _GEN_1168 : tag_143; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4776 = _T_7 ? _GEN_1169 : tag_144; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4777 = _T_7 ? _GEN_1170 : tag_145; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4778 = _T_7 ? _GEN_1171 : tag_146; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4779 = _T_7 ? _GEN_1172 : tag_147; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4780 = _T_7 ? _GEN_1173 : tag_148; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4781 = _T_7 ? _GEN_1174 : tag_149; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4782 = _T_7 ? _GEN_1175 : tag_150; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4783 = _T_7 ? _GEN_1176 : tag_151; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4784 = _T_7 ? _GEN_1177 : tag_152; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4785 = _T_7 ? _GEN_1178 : tag_153; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4786 = _T_7 ? _GEN_1179 : tag_154; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4787 = _T_7 ? _GEN_1180 : tag_155; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4788 = _T_7 ? _GEN_1181 : tag_156; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4789 = _T_7 ? _GEN_1182 : tag_157; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4790 = _T_7 ? _GEN_1183 : tag_158; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4791 = _T_7 ? _GEN_1184 : tag_159; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4792 = _T_7 ? _GEN_1185 : tag_160; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4793 = _T_7 ? _GEN_1186 : tag_161; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4794 = _T_7 ? _GEN_1187 : tag_162; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4795 = _T_7 ? _GEN_1188 : tag_163; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4796 = _T_7 ? _GEN_1189 : tag_164; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4797 = _T_7 ? _GEN_1190 : tag_165; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4798 = _T_7 ? _GEN_1191 : tag_166; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4799 = _T_7 ? _GEN_1192 : tag_167; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4800 = _T_7 ? _GEN_1193 : tag_168; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4801 = _T_7 ? _GEN_1194 : tag_169; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4802 = _T_7 ? _GEN_1195 : tag_170; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4803 = _T_7 ? _GEN_1196 : tag_171; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4804 = _T_7 ? _GEN_1197 : tag_172; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4805 = _T_7 ? _GEN_1198 : tag_173; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4806 = _T_7 ? _GEN_1199 : tag_174; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4807 = _T_7 ? _GEN_1200 : tag_175; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4808 = _T_7 ? _GEN_1201 : tag_176; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4809 = _T_7 ? _GEN_1202 : tag_177; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4810 = _T_7 ? _GEN_1203 : tag_178; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4811 = _T_7 ? _GEN_1204 : tag_179; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4812 = _T_7 ? _GEN_1205 : tag_180; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4813 = _T_7 ? _GEN_1206 : tag_181; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4814 = _T_7 ? _GEN_1207 : tag_182; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4815 = _T_7 ? _GEN_1208 : tag_183; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4816 = _T_7 ? _GEN_1209 : tag_184; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4817 = _T_7 ? _GEN_1210 : tag_185; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4818 = _T_7 ? _GEN_1211 : tag_186; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4819 = _T_7 ? _GEN_1212 : tag_187; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4820 = _T_7 ? _GEN_1213 : tag_188; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4821 = _T_7 ? _GEN_1214 : tag_189; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4822 = _T_7 ? _GEN_1215 : tag_190; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4823 = _T_7 ? _GEN_1216 : tag_191; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4824 = _T_7 ? _GEN_1217 : tag_192; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4825 = _T_7 ? _GEN_1218 : tag_193; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4826 = _T_7 ? _GEN_1219 : tag_194; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4827 = _T_7 ? _GEN_1220 : tag_195; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4828 = _T_7 ? _GEN_1221 : tag_196; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4829 = _T_7 ? _GEN_1222 : tag_197; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4830 = _T_7 ? _GEN_1223 : tag_198; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4831 = _T_7 ? _GEN_1224 : tag_199; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4832 = _T_7 ? _GEN_1225 : tag_200; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4833 = _T_7 ? _GEN_1226 : tag_201; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4834 = _T_7 ? _GEN_1227 : tag_202; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4835 = _T_7 ? _GEN_1228 : tag_203; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4836 = _T_7 ? _GEN_1229 : tag_204; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4837 = _T_7 ? _GEN_1230 : tag_205; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4838 = _T_7 ? _GEN_1231 : tag_206; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4839 = _T_7 ? _GEN_1232 : tag_207; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4840 = _T_7 ? _GEN_1233 : tag_208; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4841 = _T_7 ? _GEN_1234 : tag_209; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4842 = _T_7 ? _GEN_1235 : tag_210; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4843 = _T_7 ? _GEN_1236 : tag_211; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4844 = _T_7 ? _GEN_1237 : tag_212; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4845 = _T_7 ? _GEN_1238 : tag_213; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4846 = _T_7 ? _GEN_1239 : tag_214; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4847 = _T_7 ? _GEN_1240 : tag_215; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4848 = _T_7 ? _GEN_1241 : tag_216; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4849 = _T_7 ? _GEN_1242 : tag_217; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4850 = _T_7 ? _GEN_1243 : tag_218; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4851 = _T_7 ? _GEN_1244 : tag_219; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4852 = _T_7 ? _GEN_1245 : tag_220; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4853 = _T_7 ? _GEN_1246 : tag_221; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4854 = _T_7 ? _GEN_1247 : tag_222; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4855 = _T_7 ? _GEN_1248 : tag_223; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4856 = _T_7 ? _GEN_1249 : tag_224; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4857 = _T_7 ? _GEN_1250 : tag_225; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4858 = _T_7 ? _GEN_1251 : tag_226; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4859 = _T_7 ? _GEN_1252 : tag_227; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4860 = _T_7 ? _GEN_1253 : tag_228; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4861 = _T_7 ? _GEN_1254 : tag_229; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4862 = _T_7 ? _GEN_1255 : tag_230; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4863 = _T_7 ? _GEN_1256 : tag_231; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4864 = _T_7 ? _GEN_1257 : tag_232; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4865 = _T_7 ? _GEN_1258 : tag_233; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4866 = _T_7 ? _GEN_1259 : tag_234; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4867 = _T_7 ? _GEN_1260 : tag_235; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4868 = _T_7 ? _GEN_1261 : tag_236; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4869 = _T_7 ? _GEN_1262 : tag_237; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4870 = _T_7 ? _GEN_1263 : tag_238; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4871 = _T_7 ? _GEN_1264 : tag_239; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4872 = _T_7 ? _GEN_1265 : tag_240; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4873 = _T_7 ? _GEN_1266 : tag_241; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4874 = _T_7 ? _GEN_1267 : tag_242; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4875 = _T_7 ? _GEN_1268 : tag_243; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4876 = _T_7 ? _GEN_1269 : tag_244; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4877 = _T_7 ? _GEN_1270 : tag_245; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4878 = _T_7 ? _GEN_1271 : tag_246; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4879 = _T_7 ? _GEN_1272 : tag_247; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4880 = _T_7 ? _GEN_1273 : tag_248; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4881 = _T_7 ? _GEN_1274 : tag_249; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4882 = _T_7 ? _GEN_1275 : tag_250; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4883 = _T_7 ? _GEN_1276 : tag_251; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4884 = _T_7 ? _GEN_1277 : tag_252; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4885 = _T_7 ? _GEN_1278 : tag_253; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4886 = _T_7 ? _GEN_1279 : tag_254; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_4887 = _T_7 ? _GEN_1280 : tag_255; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire  _GEN_4888 = _T_7 ? _GEN_1537 : dirty_0; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4889 = _T_7 ? _GEN_1538 : dirty_1; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4890 = _T_7 ? _GEN_1539 : dirty_2; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4891 = _T_7 ? _GEN_1540 : dirty_3; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4892 = _T_7 ? _GEN_1541 : dirty_4; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4893 = _T_7 ? _GEN_1542 : dirty_5; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4894 = _T_7 ? _GEN_1543 : dirty_6; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4895 = _T_7 ? _GEN_1544 : dirty_7; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4896 = _T_7 ? _GEN_1545 : dirty_8; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4897 = _T_7 ? _GEN_1546 : dirty_9; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4898 = _T_7 ? _GEN_1547 : dirty_10; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4899 = _T_7 ? _GEN_1548 : dirty_11; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4900 = _T_7 ? _GEN_1549 : dirty_12; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4901 = _T_7 ? _GEN_1550 : dirty_13; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4902 = _T_7 ? _GEN_1551 : dirty_14; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4903 = _T_7 ? _GEN_1552 : dirty_15; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4904 = _T_7 ? _GEN_1553 : dirty_16; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4905 = _T_7 ? _GEN_1554 : dirty_17; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4906 = _T_7 ? _GEN_1555 : dirty_18; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4907 = _T_7 ? _GEN_1556 : dirty_19; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4908 = _T_7 ? _GEN_1557 : dirty_20; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4909 = _T_7 ? _GEN_1558 : dirty_21; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4910 = _T_7 ? _GEN_1559 : dirty_22; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4911 = _T_7 ? _GEN_1560 : dirty_23; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4912 = _T_7 ? _GEN_1561 : dirty_24; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4913 = _T_7 ? _GEN_1562 : dirty_25; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4914 = _T_7 ? _GEN_1563 : dirty_26; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4915 = _T_7 ? _GEN_1564 : dirty_27; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4916 = _T_7 ? _GEN_1565 : dirty_28; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4917 = _T_7 ? _GEN_1566 : dirty_29; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4918 = _T_7 ? _GEN_1567 : dirty_30; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4919 = _T_7 ? _GEN_1568 : dirty_31; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4920 = _T_7 ? _GEN_1569 : dirty_32; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4921 = _T_7 ? _GEN_1570 : dirty_33; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4922 = _T_7 ? _GEN_1571 : dirty_34; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4923 = _T_7 ? _GEN_1572 : dirty_35; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4924 = _T_7 ? _GEN_1573 : dirty_36; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4925 = _T_7 ? _GEN_1574 : dirty_37; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4926 = _T_7 ? _GEN_1575 : dirty_38; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4927 = _T_7 ? _GEN_1576 : dirty_39; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4928 = _T_7 ? _GEN_1577 : dirty_40; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4929 = _T_7 ? _GEN_1578 : dirty_41; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4930 = _T_7 ? _GEN_1579 : dirty_42; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4931 = _T_7 ? _GEN_1580 : dirty_43; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4932 = _T_7 ? _GEN_1581 : dirty_44; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4933 = _T_7 ? _GEN_1582 : dirty_45; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4934 = _T_7 ? _GEN_1583 : dirty_46; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4935 = _T_7 ? _GEN_1584 : dirty_47; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4936 = _T_7 ? _GEN_1585 : dirty_48; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4937 = _T_7 ? _GEN_1586 : dirty_49; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4938 = _T_7 ? _GEN_1587 : dirty_50; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4939 = _T_7 ? _GEN_1588 : dirty_51; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4940 = _T_7 ? _GEN_1589 : dirty_52; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4941 = _T_7 ? _GEN_1590 : dirty_53; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4942 = _T_7 ? _GEN_1591 : dirty_54; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4943 = _T_7 ? _GEN_1592 : dirty_55; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4944 = _T_7 ? _GEN_1593 : dirty_56; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4945 = _T_7 ? _GEN_1594 : dirty_57; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4946 = _T_7 ? _GEN_1595 : dirty_58; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4947 = _T_7 ? _GEN_1596 : dirty_59; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4948 = _T_7 ? _GEN_1597 : dirty_60; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4949 = _T_7 ? _GEN_1598 : dirty_61; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4950 = _T_7 ? _GEN_1599 : dirty_62; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4951 = _T_7 ? _GEN_1600 : dirty_63; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4952 = _T_7 ? _GEN_1601 : dirty_64; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4953 = _T_7 ? _GEN_1602 : dirty_65; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4954 = _T_7 ? _GEN_1603 : dirty_66; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4955 = _T_7 ? _GEN_1604 : dirty_67; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4956 = _T_7 ? _GEN_1605 : dirty_68; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4957 = _T_7 ? _GEN_1606 : dirty_69; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4958 = _T_7 ? _GEN_1607 : dirty_70; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4959 = _T_7 ? _GEN_1608 : dirty_71; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4960 = _T_7 ? _GEN_1609 : dirty_72; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4961 = _T_7 ? _GEN_1610 : dirty_73; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4962 = _T_7 ? _GEN_1611 : dirty_74; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4963 = _T_7 ? _GEN_1612 : dirty_75; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4964 = _T_7 ? _GEN_1613 : dirty_76; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4965 = _T_7 ? _GEN_1614 : dirty_77; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4966 = _T_7 ? _GEN_1615 : dirty_78; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4967 = _T_7 ? _GEN_1616 : dirty_79; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4968 = _T_7 ? _GEN_1617 : dirty_80; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4969 = _T_7 ? _GEN_1618 : dirty_81; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4970 = _T_7 ? _GEN_1619 : dirty_82; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4971 = _T_7 ? _GEN_1620 : dirty_83; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4972 = _T_7 ? _GEN_1621 : dirty_84; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4973 = _T_7 ? _GEN_1622 : dirty_85; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4974 = _T_7 ? _GEN_1623 : dirty_86; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4975 = _T_7 ? _GEN_1624 : dirty_87; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4976 = _T_7 ? _GEN_1625 : dirty_88; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4977 = _T_7 ? _GEN_1626 : dirty_89; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4978 = _T_7 ? _GEN_1627 : dirty_90; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4979 = _T_7 ? _GEN_1628 : dirty_91; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4980 = _T_7 ? _GEN_1629 : dirty_92; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4981 = _T_7 ? _GEN_1630 : dirty_93; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4982 = _T_7 ? _GEN_1631 : dirty_94; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4983 = _T_7 ? _GEN_1632 : dirty_95; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4984 = _T_7 ? _GEN_1633 : dirty_96; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4985 = _T_7 ? _GEN_1634 : dirty_97; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4986 = _T_7 ? _GEN_1635 : dirty_98; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4987 = _T_7 ? _GEN_1636 : dirty_99; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4988 = _T_7 ? _GEN_1637 : dirty_100; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4989 = _T_7 ? _GEN_1638 : dirty_101; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4990 = _T_7 ? _GEN_1639 : dirty_102; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4991 = _T_7 ? _GEN_1640 : dirty_103; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4992 = _T_7 ? _GEN_1641 : dirty_104; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4993 = _T_7 ? _GEN_1642 : dirty_105; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4994 = _T_7 ? _GEN_1643 : dirty_106; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4995 = _T_7 ? _GEN_1644 : dirty_107; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4996 = _T_7 ? _GEN_1645 : dirty_108; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4997 = _T_7 ? _GEN_1646 : dirty_109; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4998 = _T_7 ? _GEN_1647 : dirty_110; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_4999 = _T_7 ? _GEN_1648 : dirty_111; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5000 = _T_7 ? _GEN_1649 : dirty_112; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5001 = _T_7 ? _GEN_1650 : dirty_113; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5002 = _T_7 ? _GEN_1651 : dirty_114; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5003 = _T_7 ? _GEN_1652 : dirty_115; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5004 = _T_7 ? _GEN_1653 : dirty_116; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5005 = _T_7 ? _GEN_1654 : dirty_117; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5006 = _T_7 ? _GEN_1655 : dirty_118; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5007 = _T_7 ? _GEN_1656 : dirty_119; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5008 = _T_7 ? _GEN_1657 : dirty_120; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5009 = _T_7 ? _GEN_1658 : dirty_121; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5010 = _T_7 ? _GEN_1659 : dirty_122; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5011 = _T_7 ? _GEN_1660 : dirty_123; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5012 = _T_7 ? _GEN_1661 : dirty_124; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5013 = _T_7 ? _GEN_1662 : dirty_125; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5014 = _T_7 ? _GEN_1663 : dirty_126; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5015 = _T_7 ? _GEN_1664 : dirty_127; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5016 = _T_7 ? _GEN_1665 : dirty_128; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5017 = _T_7 ? _GEN_1666 : dirty_129; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5018 = _T_7 ? _GEN_1667 : dirty_130; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5019 = _T_7 ? _GEN_1668 : dirty_131; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5020 = _T_7 ? _GEN_1669 : dirty_132; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5021 = _T_7 ? _GEN_1670 : dirty_133; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5022 = _T_7 ? _GEN_1671 : dirty_134; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5023 = _T_7 ? _GEN_1672 : dirty_135; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5024 = _T_7 ? _GEN_1673 : dirty_136; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5025 = _T_7 ? _GEN_1674 : dirty_137; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5026 = _T_7 ? _GEN_1675 : dirty_138; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5027 = _T_7 ? _GEN_1676 : dirty_139; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5028 = _T_7 ? _GEN_1677 : dirty_140; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5029 = _T_7 ? _GEN_1678 : dirty_141; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5030 = _T_7 ? _GEN_1679 : dirty_142; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5031 = _T_7 ? _GEN_1680 : dirty_143; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5032 = _T_7 ? _GEN_1681 : dirty_144; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5033 = _T_7 ? _GEN_1682 : dirty_145; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5034 = _T_7 ? _GEN_1683 : dirty_146; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5035 = _T_7 ? _GEN_1684 : dirty_147; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5036 = _T_7 ? _GEN_1685 : dirty_148; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5037 = _T_7 ? _GEN_1686 : dirty_149; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5038 = _T_7 ? _GEN_1687 : dirty_150; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5039 = _T_7 ? _GEN_1688 : dirty_151; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5040 = _T_7 ? _GEN_1689 : dirty_152; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5041 = _T_7 ? _GEN_1690 : dirty_153; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5042 = _T_7 ? _GEN_1691 : dirty_154; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5043 = _T_7 ? _GEN_1692 : dirty_155; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5044 = _T_7 ? _GEN_1693 : dirty_156; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5045 = _T_7 ? _GEN_1694 : dirty_157; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5046 = _T_7 ? _GEN_1695 : dirty_158; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5047 = _T_7 ? _GEN_1696 : dirty_159; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5048 = _T_7 ? _GEN_1697 : dirty_160; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5049 = _T_7 ? _GEN_1698 : dirty_161; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5050 = _T_7 ? _GEN_1699 : dirty_162; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5051 = _T_7 ? _GEN_1700 : dirty_163; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5052 = _T_7 ? _GEN_1701 : dirty_164; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5053 = _T_7 ? _GEN_1702 : dirty_165; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5054 = _T_7 ? _GEN_1703 : dirty_166; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5055 = _T_7 ? _GEN_1704 : dirty_167; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5056 = _T_7 ? _GEN_1705 : dirty_168; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5057 = _T_7 ? _GEN_1706 : dirty_169; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5058 = _T_7 ? _GEN_1707 : dirty_170; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5059 = _T_7 ? _GEN_1708 : dirty_171; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5060 = _T_7 ? _GEN_1709 : dirty_172; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5061 = _T_7 ? _GEN_1710 : dirty_173; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5062 = _T_7 ? _GEN_1711 : dirty_174; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5063 = _T_7 ? _GEN_1712 : dirty_175; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5064 = _T_7 ? _GEN_1713 : dirty_176; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5065 = _T_7 ? _GEN_1714 : dirty_177; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5066 = _T_7 ? _GEN_1715 : dirty_178; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5067 = _T_7 ? _GEN_1716 : dirty_179; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5068 = _T_7 ? _GEN_1717 : dirty_180; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5069 = _T_7 ? _GEN_1718 : dirty_181; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5070 = _T_7 ? _GEN_1719 : dirty_182; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5071 = _T_7 ? _GEN_1720 : dirty_183; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5072 = _T_7 ? _GEN_1721 : dirty_184; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5073 = _T_7 ? _GEN_1722 : dirty_185; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5074 = _T_7 ? _GEN_1723 : dirty_186; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5075 = _T_7 ? _GEN_1724 : dirty_187; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5076 = _T_7 ? _GEN_1725 : dirty_188; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5077 = _T_7 ? _GEN_1726 : dirty_189; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5078 = _T_7 ? _GEN_1727 : dirty_190; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5079 = _T_7 ? _GEN_1728 : dirty_191; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5080 = _T_7 ? _GEN_1729 : dirty_192; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5081 = _T_7 ? _GEN_1730 : dirty_193; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5082 = _T_7 ? _GEN_1731 : dirty_194; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5083 = _T_7 ? _GEN_1732 : dirty_195; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5084 = _T_7 ? _GEN_1733 : dirty_196; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5085 = _T_7 ? _GEN_1734 : dirty_197; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5086 = _T_7 ? _GEN_1735 : dirty_198; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5087 = _T_7 ? _GEN_1736 : dirty_199; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5088 = _T_7 ? _GEN_1737 : dirty_200; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5089 = _T_7 ? _GEN_1738 : dirty_201; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5090 = _T_7 ? _GEN_1739 : dirty_202; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5091 = _T_7 ? _GEN_1740 : dirty_203; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5092 = _T_7 ? _GEN_1741 : dirty_204; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5093 = _T_7 ? _GEN_1742 : dirty_205; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5094 = _T_7 ? _GEN_1743 : dirty_206; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5095 = _T_7 ? _GEN_1744 : dirty_207; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5096 = _T_7 ? _GEN_1745 : dirty_208; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5097 = _T_7 ? _GEN_1746 : dirty_209; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5098 = _T_7 ? _GEN_1747 : dirty_210; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5099 = _T_7 ? _GEN_1748 : dirty_211; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5100 = _T_7 ? _GEN_1749 : dirty_212; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5101 = _T_7 ? _GEN_1750 : dirty_213; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5102 = _T_7 ? _GEN_1751 : dirty_214; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5103 = _T_7 ? _GEN_1752 : dirty_215; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5104 = _T_7 ? _GEN_1753 : dirty_216; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5105 = _T_7 ? _GEN_1754 : dirty_217; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5106 = _T_7 ? _GEN_1755 : dirty_218; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5107 = _T_7 ? _GEN_1756 : dirty_219; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5108 = _T_7 ? _GEN_1757 : dirty_220; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5109 = _T_7 ? _GEN_1758 : dirty_221; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5110 = _T_7 ? _GEN_1759 : dirty_222; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5111 = _T_7 ? _GEN_1760 : dirty_223; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5112 = _T_7 ? _GEN_1761 : dirty_224; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5113 = _T_7 ? _GEN_1762 : dirty_225; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5114 = _T_7 ? _GEN_1763 : dirty_226; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5115 = _T_7 ? _GEN_1764 : dirty_227; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5116 = _T_7 ? _GEN_1765 : dirty_228; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5117 = _T_7 ? _GEN_1766 : dirty_229; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5118 = _T_7 ? _GEN_1767 : dirty_230; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5119 = _T_7 ? _GEN_1768 : dirty_231; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5120 = _T_7 ? _GEN_1769 : dirty_232; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5121 = _T_7 ? _GEN_1770 : dirty_233; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5122 = _T_7 ? _GEN_1771 : dirty_234; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5123 = _T_7 ? _GEN_1772 : dirty_235; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5124 = _T_7 ? _GEN_1773 : dirty_236; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5125 = _T_7 ? _GEN_1774 : dirty_237; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5126 = _T_7 ? _GEN_1775 : dirty_238; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5127 = _T_7 ? _GEN_1776 : dirty_239; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5128 = _T_7 ? _GEN_1777 : dirty_240; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5129 = _T_7 ? _GEN_1778 : dirty_241; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5130 = _T_7 ? _GEN_1779 : dirty_242; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5131 = _T_7 ? _GEN_1780 : dirty_243; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5132 = _T_7 ? _GEN_1781 : dirty_244; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5133 = _T_7 ? _GEN_1782 : dirty_245; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5134 = _T_7 ? _GEN_1783 : dirty_246; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5135 = _T_7 ? _GEN_1784 : dirty_247; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5136 = _T_7 ? _GEN_1785 : dirty_248; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5137 = _T_7 ? _GEN_1786 : dirty_249; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5138 = _T_7 ? _GEN_1787 : dirty_250; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5139 = _T_7 ? _GEN_1788 : dirty_251; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5140 = _T_7 ? _GEN_1789 : dirty_252; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5141 = _T_7 ? _GEN_1790 : dirty_253; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5142 = _T_7 ? _GEN_1791 : dirty_254; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5143 = _T_7 ? _GEN_1792 : dirty_255; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire [3:0] _GEN_5144 = _T_7 ? _GEN_1281 : offset_0; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5145 = _T_7 ? _GEN_1282 : offset_1; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5146 = _T_7 ? _GEN_1283 : offset_2; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5147 = _T_7 ? _GEN_1284 : offset_3; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5148 = _T_7 ? _GEN_1285 : offset_4; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5149 = _T_7 ? _GEN_1286 : offset_5; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5150 = _T_7 ? _GEN_1287 : offset_6; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5151 = _T_7 ? _GEN_1288 : offset_7; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5152 = _T_7 ? _GEN_1289 : offset_8; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5153 = _T_7 ? _GEN_1290 : offset_9; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5154 = _T_7 ? _GEN_1291 : offset_10; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5155 = _T_7 ? _GEN_1292 : offset_11; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5156 = _T_7 ? _GEN_1293 : offset_12; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5157 = _T_7 ? _GEN_1294 : offset_13; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5158 = _T_7 ? _GEN_1295 : offset_14; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5159 = _T_7 ? _GEN_1296 : offset_15; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5160 = _T_7 ? _GEN_1297 : offset_16; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5161 = _T_7 ? _GEN_1298 : offset_17; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5162 = _T_7 ? _GEN_1299 : offset_18; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5163 = _T_7 ? _GEN_1300 : offset_19; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5164 = _T_7 ? _GEN_1301 : offset_20; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5165 = _T_7 ? _GEN_1302 : offset_21; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5166 = _T_7 ? _GEN_1303 : offset_22; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5167 = _T_7 ? _GEN_1304 : offset_23; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5168 = _T_7 ? _GEN_1305 : offset_24; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5169 = _T_7 ? _GEN_1306 : offset_25; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5170 = _T_7 ? _GEN_1307 : offset_26; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5171 = _T_7 ? _GEN_1308 : offset_27; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5172 = _T_7 ? _GEN_1309 : offset_28; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5173 = _T_7 ? _GEN_1310 : offset_29; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5174 = _T_7 ? _GEN_1311 : offset_30; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5175 = _T_7 ? _GEN_1312 : offset_31; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5176 = _T_7 ? _GEN_1313 : offset_32; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5177 = _T_7 ? _GEN_1314 : offset_33; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5178 = _T_7 ? _GEN_1315 : offset_34; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5179 = _T_7 ? _GEN_1316 : offset_35; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5180 = _T_7 ? _GEN_1317 : offset_36; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5181 = _T_7 ? _GEN_1318 : offset_37; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5182 = _T_7 ? _GEN_1319 : offset_38; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5183 = _T_7 ? _GEN_1320 : offset_39; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5184 = _T_7 ? _GEN_1321 : offset_40; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5185 = _T_7 ? _GEN_1322 : offset_41; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5186 = _T_7 ? _GEN_1323 : offset_42; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5187 = _T_7 ? _GEN_1324 : offset_43; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5188 = _T_7 ? _GEN_1325 : offset_44; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5189 = _T_7 ? _GEN_1326 : offset_45; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5190 = _T_7 ? _GEN_1327 : offset_46; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5191 = _T_7 ? _GEN_1328 : offset_47; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5192 = _T_7 ? _GEN_1329 : offset_48; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5193 = _T_7 ? _GEN_1330 : offset_49; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5194 = _T_7 ? _GEN_1331 : offset_50; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5195 = _T_7 ? _GEN_1332 : offset_51; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5196 = _T_7 ? _GEN_1333 : offset_52; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5197 = _T_7 ? _GEN_1334 : offset_53; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5198 = _T_7 ? _GEN_1335 : offset_54; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5199 = _T_7 ? _GEN_1336 : offset_55; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5200 = _T_7 ? _GEN_1337 : offset_56; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5201 = _T_7 ? _GEN_1338 : offset_57; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5202 = _T_7 ? _GEN_1339 : offset_58; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5203 = _T_7 ? _GEN_1340 : offset_59; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5204 = _T_7 ? _GEN_1341 : offset_60; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5205 = _T_7 ? _GEN_1342 : offset_61; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5206 = _T_7 ? _GEN_1343 : offset_62; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5207 = _T_7 ? _GEN_1344 : offset_63; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5208 = _T_7 ? _GEN_1345 : offset_64; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5209 = _T_7 ? _GEN_1346 : offset_65; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5210 = _T_7 ? _GEN_1347 : offset_66; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5211 = _T_7 ? _GEN_1348 : offset_67; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5212 = _T_7 ? _GEN_1349 : offset_68; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5213 = _T_7 ? _GEN_1350 : offset_69; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5214 = _T_7 ? _GEN_1351 : offset_70; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5215 = _T_7 ? _GEN_1352 : offset_71; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5216 = _T_7 ? _GEN_1353 : offset_72; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5217 = _T_7 ? _GEN_1354 : offset_73; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5218 = _T_7 ? _GEN_1355 : offset_74; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5219 = _T_7 ? _GEN_1356 : offset_75; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5220 = _T_7 ? _GEN_1357 : offset_76; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5221 = _T_7 ? _GEN_1358 : offset_77; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5222 = _T_7 ? _GEN_1359 : offset_78; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5223 = _T_7 ? _GEN_1360 : offset_79; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5224 = _T_7 ? _GEN_1361 : offset_80; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5225 = _T_7 ? _GEN_1362 : offset_81; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5226 = _T_7 ? _GEN_1363 : offset_82; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5227 = _T_7 ? _GEN_1364 : offset_83; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5228 = _T_7 ? _GEN_1365 : offset_84; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5229 = _T_7 ? _GEN_1366 : offset_85; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5230 = _T_7 ? _GEN_1367 : offset_86; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5231 = _T_7 ? _GEN_1368 : offset_87; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5232 = _T_7 ? _GEN_1369 : offset_88; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5233 = _T_7 ? _GEN_1370 : offset_89; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5234 = _T_7 ? _GEN_1371 : offset_90; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5235 = _T_7 ? _GEN_1372 : offset_91; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5236 = _T_7 ? _GEN_1373 : offset_92; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5237 = _T_7 ? _GEN_1374 : offset_93; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5238 = _T_7 ? _GEN_1375 : offset_94; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5239 = _T_7 ? _GEN_1376 : offset_95; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5240 = _T_7 ? _GEN_1377 : offset_96; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5241 = _T_7 ? _GEN_1378 : offset_97; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5242 = _T_7 ? _GEN_1379 : offset_98; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5243 = _T_7 ? _GEN_1380 : offset_99; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5244 = _T_7 ? _GEN_1381 : offset_100; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5245 = _T_7 ? _GEN_1382 : offset_101; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5246 = _T_7 ? _GEN_1383 : offset_102; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5247 = _T_7 ? _GEN_1384 : offset_103; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5248 = _T_7 ? _GEN_1385 : offset_104; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5249 = _T_7 ? _GEN_1386 : offset_105; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5250 = _T_7 ? _GEN_1387 : offset_106; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5251 = _T_7 ? _GEN_1388 : offset_107; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5252 = _T_7 ? _GEN_1389 : offset_108; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5253 = _T_7 ? _GEN_1390 : offset_109; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5254 = _T_7 ? _GEN_1391 : offset_110; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5255 = _T_7 ? _GEN_1392 : offset_111; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5256 = _T_7 ? _GEN_1393 : offset_112; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5257 = _T_7 ? _GEN_1394 : offset_113; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5258 = _T_7 ? _GEN_1395 : offset_114; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5259 = _T_7 ? _GEN_1396 : offset_115; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5260 = _T_7 ? _GEN_1397 : offset_116; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5261 = _T_7 ? _GEN_1398 : offset_117; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5262 = _T_7 ? _GEN_1399 : offset_118; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5263 = _T_7 ? _GEN_1400 : offset_119; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5264 = _T_7 ? _GEN_1401 : offset_120; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5265 = _T_7 ? _GEN_1402 : offset_121; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5266 = _T_7 ? _GEN_1403 : offset_122; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5267 = _T_7 ? _GEN_1404 : offset_123; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5268 = _T_7 ? _GEN_1405 : offset_124; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5269 = _T_7 ? _GEN_1406 : offset_125; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5270 = _T_7 ? _GEN_1407 : offset_126; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5271 = _T_7 ? _GEN_1408 : offset_127; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5272 = _T_7 ? _GEN_1409 : offset_128; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5273 = _T_7 ? _GEN_1410 : offset_129; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5274 = _T_7 ? _GEN_1411 : offset_130; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5275 = _T_7 ? _GEN_1412 : offset_131; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5276 = _T_7 ? _GEN_1413 : offset_132; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5277 = _T_7 ? _GEN_1414 : offset_133; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5278 = _T_7 ? _GEN_1415 : offset_134; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5279 = _T_7 ? _GEN_1416 : offset_135; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5280 = _T_7 ? _GEN_1417 : offset_136; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5281 = _T_7 ? _GEN_1418 : offset_137; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5282 = _T_7 ? _GEN_1419 : offset_138; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5283 = _T_7 ? _GEN_1420 : offset_139; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5284 = _T_7 ? _GEN_1421 : offset_140; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5285 = _T_7 ? _GEN_1422 : offset_141; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5286 = _T_7 ? _GEN_1423 : offset_142; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5287 = _T_7 ? _GEN_1424 : offset_143; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5288 = _T_7 ? _GEN_1425 : offset_144; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5289 = _T_7 ? _GEN_1426 : offset_145; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5290 = _T_7 ? _GEN_1427 : offset_146; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5291 = _T_7 ? _GEN_1428 : offset_147; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5292 = _T_7 ? _GEN_1429 : offset_148; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5293 = _T_7 ? _GEN_1430 : offset_149; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5294 = _T_7 ? _GEN_1431 : offset_150; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5295 = _T_7 ? _GEN_1432 : offset_151; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5296 = _T_7 ? _GEN_1433 : offset_152; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5297 = _T_7 ? _GEN_1434 : offset_153; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5298 = _T_7 ? _GEN_1435 : offset_154; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5299 = _T_7 ? _GEN_1436 : offset_155; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5300 = _T_7 ? _GEN_1437 : offset_156; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5301 = _T_7 ? _GEN_1438 : offset_157; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5302 = _T_7 ? _GEN_1439 : offset_158; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5303 = _T_7 ? _GEN_1440 : offset_159; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5304 = _T_7 ? _GEN_1441 : offset_160; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5305 = _T_7 ? _GEN_1442 : offset_161; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5306 = _T_7 ? _GEN_1443 : offset_162; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5307 = _T_7 ? _GEN_1444 : offset_163; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5308 = _T_7 ? _GEN_1445 : offset_164; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5309 = _T_7 ? _GEN_1446 : offset_165; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5310 = _T_7 ? _GEN_1447 : offset_166; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5311 = _T_7 ? _GEN_1448 : offset_167; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5312 = _T_7 ? _GEN_1449 : offset_168; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5313 = _T_7 ? _GEN_1450 : offset_169; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5314 = _T_7 ? _GEN_1451 : offset_170; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5315 = _T_7 ? _GEN_1452 : offset_171; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5316 = _T_7 ? _GEN_1453 : offset_172; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5317 = _T_7 ? _GEN_1454 : offset_173; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5318 = _T_7 ? _GEN_1455 : offset_174; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5319 = _T_7 ? _GEN_1456 : offset_175; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5320 = _T_7 ? _GEN_1457 : offset_176; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5321 = _T_7 ? _GEN_1458 : offset_177; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5322 = _T_7 ? _GEN_1459 : offset_178; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5323 = _T_7 ? _GEN_1460 : offset_179; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5324 = _T_7 ? _GEN_1461 : offset_180; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5325 = _T_7 ? _GEN_1462 : offset_181; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5326 = _T_7 ? _GEN_1463 : offset_182; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5327 = _T_7 ? _GEN_1464 : offset_183; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5328 = _T_7 ? _GEN_1465 : offset_184; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5329 = _T_7 ? _GEN_1466 : offset_185; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5330 = _T_7 ? _GEN_1467 : offset_186; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5331 = _T_7 ? _GEN_1468 : offset_187; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5332 = _T_7 ? _GEN_1469 : offset_188; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5333 = _T_7 ? _GEN_1470 : offset_189; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5334 = _T_7 ? _GEN_1471 : offset_190; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5335 = _T_7 ? _GEN_1472 : offset_191; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5336 = _T_7 ? _GEN_1473 : offset_192; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5337 = _T_7 ? _GEN_1474 : offset_193; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5338 = _T_7 ? _GEN_1475 : offset_194; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5339 = _T_7 ? _GEN_1476 : offset_195; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5340 = _T_7 ? _GEN_1477 : offset_196; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5341 = _T_7 ? _GEN_1478 : offset_197; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5342 = _T_7 ? _GEN_1479 : offset_198; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5343 = _T_7 ? _GEN_1480 : offset_199; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5344 = _T_7 ? _GEN_1481 : offset_200; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5345 = _T_7 ? _GEN_1482 : offset_201; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5346 = _T_7 ? _GEN_1483 : offset_202; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5347 = _T_7 ? _GEN_1484 : offset_203; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5348 = _T_7 ? _GEN_1485 : offset_204; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5349 = _T_7 ? _GEN_1486 : offset_205; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5350 = _T_7 ? _GEN_1487 : offset_206; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5351 = _T_7 ? _GEN_1488 : offset_207; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5352 = _T_7 ? _GEN_1489 : offset_208; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5353 = _T_7 ? _GEN_1490 : offset_209; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5354 = _T_7 ? _GEN_1491 : offset_210; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5355 = _T_7 ? _GEN_1492 : offset_211; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5356 = _T_7 ? _GEN_1493 : offset_212; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5357 = _T_7 ? _GEN_1494 : offset_213; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5358 = _T_7 ? _GEN_1495 : offset_214; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5359 = _T_7 ? _GEN_1496 : offset_215; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5360 = _T_7 ? _GEN_1497 : offset_216; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5361 = _T_7 ? _GEN_1498 : offset_217; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5362 = _T_7 ? _GEN_1499 : offset_218; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5363 = _T_7 ? _GEN_1500 : offset_219; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5364 = _T_7 ? _GEN_1501 : offset_220; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5365 = _T_7 ? _GEN_1502 : offset_221; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5366 = _T_7 ? _GEN_1503 : offset_222; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5367 = _T_7 ? _GEN_1504 : offset_223; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5368 = _T_7 ? _GEN_1505 : offset_224; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5369 = _T_7 ? _GEN_1506 : offset_225; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5370 = _T_7 ? _GEN_1507 : offset_226; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5371 = _T_7 ? _GEN_1508 : offset_227; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5372 = _T_7 ? _GEN_1509 : offset_228; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5373 = _T_7 ? _GEN_1510 : offset_229; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5374 = _T_7 ? _GEN_1511 : offset_230; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5375 = _T_7 ? _GEN_1512 : offset_231; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5376 = _T_7 ? _GEN_1513 : offset_232; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5377 = _T_7 ? _GEN_1514 : offset_233; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5378 = _T_7 ? _GEN_1515 : offset_234; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5379 = _T_7 ? _GEN_1516 : offset_235; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5380 = _T_7 ? _GEN_1517 : offset_236; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5381 = _T_7 ? _GEN_1518 : offset_237; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5382 = _T_7 ? _GEN_1519 : offset_238; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5383 = _T_7 ? _GEN_1520 : offset_239; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5384 = _T_7 ? _GEN_1521 : offset_240; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5385 = _T_7 ? _GEN_1522 : offset_241; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5386 = _T_7 ? _GEN_1523 : offset_242; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5387 = _T_7 ? _GEN_1524 : offset_243; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5388 = _T_7 ? _GEN_1525 : offset_244; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5389 = _T_7 ? _GEN_1526 : offset_245; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5390 = _T_7 ? _GEN_1527 : offset_246; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5391 = _T_7 ? _GEN_1528 : offset_247; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5392 = _T_7 ? _GEN_1529 : offset_248; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5393 = _T_7 ? _GEN_1530 : offset_249; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5394 = _T_7 ? _GEN_1531 : offset_250; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5395 = _T_7 ? _GEN_1532 : offset_251; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5396 = _T_7 ? _GEN_1533 : offset_252; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5397 = _T_7 ? _GEN_1534 : offset_253; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5398 = _T_7 ? _GEN_1535 : offset_254; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_5399 = _T_7 ? _GEN_1536 : offset_255; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [2:0] _GEN_5400 = _T_7 ? 3'h0 : state; // @[Conditional.scala 39:67 Dcache.scala 203:25 Dcache.scala 26:22]
  wire [2:0] _GEN_5401 = _T_5 ? _GEN_3337 : _GEN_5400; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_5402 = _T_5 ? _GEN_3338 : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_5408 = _T_5 ? _GEN_3344 : _GEN_4373; // @[Conditional.scala 39:67]
  wire  _GEN_5409 = _T_5 ? _GEN_3345 : _GEN_4375; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_5410 = _T_5 ? _GEN_3346 : cache_wdata; // @[Conditional.scala 39:67 Dcache.scala 118:28]
  wire [127:0] _GEN_5411 = _T_5 ? _GEN_3347 : cache_strb; // @[Conditional.scala 39:67 Dcache.scala 119:28]
  wire  _GEN_5412 = _T_5 ? data_ready : _GEN_4374; // @[Conditional.scala 39:67 Dcache.scala 46:28]
  wire  _GEN_5413 = _T_5 ? valid_0 : _GEN_4376; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5414 = _T_5 ? valid_1 : _GEN_4377; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5415 = _T_5 ? valid_2 : _GEN_4378; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5416 = _T_5 ? valid_3 : _GEN_4379; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5417 = _T_5 ? valid_4 : _GEN_4380; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5418 = _T_5 ? valid_5 : _GEN_4381; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5419 = _T_5 ? valid_6 : _GEN_4382; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5420 = _T_5 ? valid_7 : _GEN_4383; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5421 = _T_5 ? valid_8 : _GEN_4384; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5422 = _T_5 ? valid_9 : _GEN_4385; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5423 = _T_5 ? valid_10 : _GEN_4386; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5424 = _T_5 ? valid_11 : _GEN_4387; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5425 = _T_5 ? valid_12 : _GEN_4388; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5426 = _T_5 ? valid_13 : _GEN_4389; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5427 = _T_5 ? valid_14 : _GEN_4390; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5428 = _T_5 ? valid_15 : _GEN_4391; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5429 = _T_5 ? valid_16 : _GEN_4392; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5430 = _T_5 ? valid_17 : _GEN_4393; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5431 = _T_5 ? valid_18 : _GEN_4394; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5432 = _T_5 ? valid_19 : _GEN_4395; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5433 = _T_5 ? valid_20 : _GEN_4396; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5434 = _T_5 ? valid_21 : _GEN_4397; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5435 = _T_5 ? valid_22 : _GEN_4398; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5436 = _T_5 ? valid_23 : _GEN_4399; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5437 = _T_5 ? valid_24 : _GEN_4400; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5438 = _T_5 ? valid_25 : _GEN_4401; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5439 = _T_5 ? valid_26 : _GEN_4402; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5440 = _T_5 ? valid_27 : _GEN_4403; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5441 = _T_5 ? valid_28 : _GEN_4404; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5442 = _T_5 ? valid_29 : _GEN_4405; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5443 = _T_5 ? valid_30 : _GEN_4406; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5444 = _T_5 ? valid_31 : _GEN_4407; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5445 = _T_5 ? valid_32 : _GEN_4408; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5446 = _T_5 ? valid_33 : _GEN_4409; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5447 = _T_5 ? valid_34 : _GEN_4410; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5448 = _T_5 ? valid_35 : _GEN_4411; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5449 = _T_5 ? valid_36 : _GEN_4412; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5450 = _T_5 ? valid_37 : _GEN_4413; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5451 = _T_5 ? valid_38 : _GEN_4414; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5452 = _T_5 ? valid_39 : _GEN_4415; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5453 = _T_5 ? valid_40 : _GEN_4416; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5454 = _T_5 ? valid_41 : _GEN_4417; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5455 = _T_5 ? valid_42 : _GEN_4418; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5456 = _T_5 ? valid_43 : _GEN_4419; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5457 = _T_5 ? valid_44 : _GEN_4420; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5458 = _T_5 ? valid_45 : _GEN_4421; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5459 = _T_5 ? valid_46 : _GEN_4422; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5460 = _T_5 ? valid_47 : _GEN_4423; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5461 = _T_5 ? valid_48 : _GEN_4424; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5462 = _T_5 ? valid_49 : _GEN_4425; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5463 = _T_5 ? valid_50 : _GEN_4426; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5464 = _T_5 ? valid_51 : _GEN_4427; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5465 = _T_5 ? valid_52 : _GEN_4428; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5466 = _T_5 ? valid_53 : _GEN_4429; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5467 = _T_5 ? valid_54 : _GEN_4430; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5468 = _T_5 ? valid_55 : _GEN_4431; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5469 = _T_5 ? valid_56 : _GEN_4432; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5470 = _T_5 ? valid_57 : _GEN_4433; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5471 = _T_5 ? valid_58 : _GEN_4434; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5472 = _T_5 ? valid_59 : _GEN_4435; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5473 = _T_5 ? valid_60 : _GEN_4436; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5474 = _T_5 ? valid_61 : _GEN_4437; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5475 = _T_5 ? valid_62 : _GEN_4438; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5476 = _T_5 ? valid_63 : _GEN_4439; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5477 = _T_5 ? valid_64 : _GEN_4440; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5478 = _T_5 ? valid_65 : _GEN_4441; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5479 = _T_5 ? valid_66 : _GEN_4442; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5480 = _T_5 ? valid_67 : _GEN_4443; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5481 = _T_5 ? valid_68 : _GEN_4444; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5482 = _T_5 ? valid_69 : _GEN_4445; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5483 = _T_5 ? valid_70 : _GEN_4446; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5484 = _T_5 ? valid_71 : _GEN_4447; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5485 = _T_5 ? valid_72 : _GEN_4448; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5486 = _T_5 ? valid_73 : _GEN_4449; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5487 = _T_5 ? valid_74 : _GEN_4450; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5488 = _T_5 ? valid_75 : _GEN_4451; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5489 = _T_5 ? valid_76 : _GEN_4452; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5490 = _T_5 ? valid_77 : _GEN_4453; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5491 = _T_5 ? valid_78 : _GEN_4454; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5492 = _T_5 ? valid_79 : _GEN_4455; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5493 = _T_5 ? valid_80 : _GEN_4456; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5494 = _T_5 ? valid_81 : _GEN_4457; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5495 = _T_5 ? valid_82 : _GEN_4458; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5496 = _T_5 ? valid_83 : _GEN_4459; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5497 = _T_5 ? valid_84 : _GEN_4460; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5498 = _T_5 ? valid_85 : _GEN_4461; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5499 = _T_5 ? valid_86 : _GEN_4462; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5500 = _T_5 ? valid_87 : _GEN_4463; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5501 = _T_5 ? valid_88 : _GEN_4464; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5502 = _T_5 ? valid_89 : _GEN_4465; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5503 = _T_5 ? valid_90 : _GEN_4466; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5504 = _T_5 ? valid_91 : _GEN_4467; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5505 = _T_5 ? valid_92 : _GEN_4468; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5506 = _T_5 ? valid_93 : _GEN_4469; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5507 = _T_5 ? valid_94 : _GEN_4470; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5508 = _T_5 ? valid_95 : _GEN_4471; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5509 = _T_5 ? valid_96 : _GEN_4472; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5510 = _T_5 ? valid_97 : _GEN_4473; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5511 = _T_5 ? valid_98 : _GEN_4474; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5512 = _T_5 ? valid_99 : _GEN_4475; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5513 = _T_5 ? valid_100 : _GEN_4476; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5514 = _T_5 ? valid_101 : _GEN_4477; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5515 = _T_5 ? valid_102 : _GEN_4478; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5516 = _T_5 ? valid_103 : _GEN_4479; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5517 = _T_5 ? valid_104 : _GEN_4480; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5518 = _T_5 ? valid_105 : _GEN_4481; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5519 = _T_5 ? valid_106 : _GEN_4482; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5520 = _T_5 ? valid_107 : _GEN_4483; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5521 = _T_5 ? valid_108 : _GEN_4484; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5522 = _T_5 ? valid_109 : _GEN_4485; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5523 = _T_5 ? valid_110 : _GEN_4486; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5524 = _T_5 ? valid_111 : _GEN_4487; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5525 = _T_5 ? valid_112 : _GEN_4488; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5526 = _T_5 ? valid_113 : _GEN_4489; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5527 = _T_5 ? valid_114 : _GEN_4490; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5528 = _T_5 ? valid_115 : _GEN_4491; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5529 = _T_5 ? valid_116 : _GEN_4492; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5530 = _T_5 ? valid_117 : _GEN_4493; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5531 = _T_5 ? valid_118 : _GEN_4494; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5532 = _T_5 ? valid_119 : _GEN_4495; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5533 = _T_5 ? valid_120 : _GEN_4496; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5534 = _T_5 ? valid_121 : _GEN_4497; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5535 = _T_5 ? valid_122 : _GEN_4498; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5536 = _T_5 ? valid_123 : _GEN_4499; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5537 = _T_5 ? valid_124 : _GEN_4500; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5538 = _T_5 ? valid_125 : _GEN_4501; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5539 = _T_5 ? valid_126 : _GEN_4502; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5540 = _T_5 ? valid_127 : _GEN_4503; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5541 = _T_5 ? valid_128 : _GEN_4504; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5542 = _T_5 ? valid_129 : _GEN_4505; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5543 = _T_5 ? valid_130 : _GEN_4506; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5544 = _T_5 ? valid_131 : _GEN_4507; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5545 = _T_5 ? valid_132 : _GEN_4508; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5546 = _T_5 ? valid_133 : _GEN_4509; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5547 = _T_5 ? valid_134 : _GEN_4510; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5548 = _T_5 ? valid_135 : _GEN_4511; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5549 = _T_5 ? valid_136 : _GEN_4512; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5550 = _T_5 ? valid_137 : _GEN_4513; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5551 = _T_5 ? valid_138 : _GEN_4514; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5552 = _T_5 ? valid_139 : _GEN_4515; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5553 = _T_5 ? valid_140 : _GEN_4516; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5554 = _T_5 ? valid_141 : _GEN_4517; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5555 = _T_5 ? valid_142 : _GEN_4518; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5556 = _T_5 ? valid_143 : _GEN_4519; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5557 = _T_5 ? valid_144 : _GEN_4520; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5558 = _T_5 ? valid_145 : _GEN_4521; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5559 = _T_5 ? valid_146 : _GEN_4522; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5560 = _T_5 ? valid_147 : _GEN_4523; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5561 = _T_5 ? valid_148 : _GEN_4524; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5562 = _T_5 ? valid_149 : _GEN_4525; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5563 = _T_5 ? valid_150 : _GEN_4526; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5564 = _T_5 ? valid_151 : _GEN_4527; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5565 = _T_5 ? valid_152 : _GEN_4528; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5566 = _T_5 ? valid_153 : _GEN_4529; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5567 = _T_5 ? valid_154 : _GEN_4530; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5568 = _T_5 ? valid_155 : _GEN_4531; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5569 = _T_5 ? valid_156 : _GEN_4532; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5570 = _T_5 ? valid_157 : _GEN_4533; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5571 = _T_5 ? valid_158 : _GEN_4534; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5572 = _T_5 ? valid_159 : _GEN_4535; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5573 = _T_5 ? valid_160 : _GEN_4536; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5574 = _T_5 ? valid_161 : _GEN_4537; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5575 = _T_5 ? valid_162 : _GEN_4538; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5576 = _T_5 ? valid_163 : _GEN_4539; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5577 = _T_5 ? valid_164 : _GEN_4540; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5578 = _T_5 ? valid_165 : _GEN_4541; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5579 = _T_5 ? valid_166 : _GEN_4542; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5580 = _T_5 ? valid_167 : _GEN_4543; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5581 = _T_5 ? valid_168 : _GEN_4544; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5582 = _T_5 ? valid_169 : _GEN_4545; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5583 = _T_5 ? valid_170 : _GEN_4546; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5584 = _T_5 ? valid_171 : _GEN_4547; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5585 = _T_5 ? valid_172 : _GEN_4548; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5586 = _T_5 ? valid_173 : _GEN_4549; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5587 = _T_5 ? valid_174 : _GEN_4550; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5588 = _T_5 ? valid_175 : _GEN_4551; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5589 = _T_5 ? valid_176 : _GEN_4552; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5590 = _T_5 ? valid_177 : _GEN_4553; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5591 = _T_5 ? valid_178 : _GEN_4554; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5592 = _T_5 ? valid_179 : _GEN_4555; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5593 = _T_5 ? valid_180 : _GEN_4556; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5594 = _T_5 ? valid_181 : _GEN_4557; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5595 = _T_5 ? valid_182 : _GEN_4558; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5596 = _T_5 ? valid_183 : _GEN_4559; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5597 = _T_5 ? valid_184 : _GEN_4560; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5598 = _T_5 ? valid_185 : _GEN_4561; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5599 = _T_5 ? valid_186 : _GEN_4562; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5600 = _T_5 ? valid_187 : _GEN_4563; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5601 = _T_5 ? valid_188 : _GEN_4564; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5602 = _T_5 ? valid_189 : _GEN_4565; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5603 = _T_5 ? valid_190 : _GEN_4566; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5604 = _T_5 ? valid_191 : _GEN_4567; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5605 = _T_5 ? valid_192 : _GEN_4568; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5606 = _T_5 ? valid_193 : _GEN_4569; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5607 = _T_5 ? valid_194 : _GEN_4570; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5608 = _T_5 ? valid_195 : _GEN_4571; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5609 = _T_5 ? valid_196 : _GEN_4572; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5610 = _T_5 ? valid_197 : _GEN_4573; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5611 = _T_5 ? valid_198 : _GEN_4574; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5612 = _T_5 ? valid_199 : _GEN_4575; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5613 = _T_5 ? valid_200 : _GEN_4576; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5614 = _T_5 ? valid_201 : _GEN_4577; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5615 = _T_5 ? valid_202 : _GEN_4578; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5616 = _T_5 ? valid_203 : _GEN_4579; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5617 = _T_5 ? valid_204 : _GEN_4580; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5618 = _T_5 ? valid_205 : _GEN_4581; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5619 = _T_5 ? valid_206 : _GEN_4582; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5620 = _T_5 ? valid_207 : _GEN_4583; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5621 = _T_5 ? valid_208 : _GEN_4584; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5622 = _T_5 ? valid_209 : _GEN_4585; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5623 = _T_5 ? valid_210 : _GEN_4586; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5624 = _T_5 ? valid_211 : _GEN_4587; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5625 = _T_5 ? valid_212 : _GEN_4588; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5626 = _T_5 ? valid_213 : _GEN_4589; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5627 = _T_5 ? valid_214 : _GEN_4590; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5628 = _T_5 ? valid_215 : _GEN_4591; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5629 = _T_5 ? valid_216 : _GEN_4592; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5630 = _T_5 ? valid_217 : _GEN_4593; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5631 = _T_5 ? valid_218 : _GEN_4594; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5632 = _T_5 ? valid_219 : _GEN_4595; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5633 = _T_5 ? valid_220 : _GEN_4596; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5634 = _T_5 ? valid_221 : _GEN_4597; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5635 = _T_5 ? valid_222 : _GEN_4598; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5636 = _T_5 ? valid_223 : _GEN_4599; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5637 = _T_5 ? valid_224 : _GEN_4600; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5638 = _T_5 ? valid_225 : _GEN_4601; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5639 = _T_5 ? valid_226 : _GEN_4602; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5640 = _T_5 ? valid_227 : _GEN_4603; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5641 = _T_5 ? valid_228 : _GEN_4604; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5642 = _T_5 ? valid_229 : _GEN_4605; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5643 = _T_5 ? valid_230 : _GEN_4606; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5644 = _T_5 ? valid_231 : _GEN_4607; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5645 = _T_5 ? valid_232 : _GEN_4608; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5646 = _T_5 ? valid_233 : _GEN_4609; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5647 = _T_5 ? valid_234 : _GEN_4610; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5648 = _T_5 ? valid_235 : _GEN_4611; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5649 = _T_5 ? valid_236 : _GEN_4612; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5650 = _T_5 ? valid_237 : _GEN_4613; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5651 = _T_5 ? valid_238 : _GEN_4614; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5652 = _T_5 ? valid_239 : _GEN_4615; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5653 = _T_5 ? valid_240 : _GEN_4616; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5654 = _T_5 ? valid_241 : _GEN_4617; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5655 = _T_5 ? valid_242 : _GEN_4618; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5656 = _T_5 ? valid_243 : _GEN_4619; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5657 = _T_5 ? valid_244 : _GEN_4620; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5658 = _T_5 ? valid_245 : _GEN_4621; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5659 = _T_5 ? valid_246 : _GEN_4622; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5660 = _T_5 ? valid_247 : _GEN_4623; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5661 = _T_5 ? valid_248 : _GEN_4624; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5662 = _T_5 ? valid_249 : _GEN_4625; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5663 = _T_5 ? valid_250 : _GEN_4626; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5664 = _T_5 ? valid_251 : _GEN_4627; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5665 = _T_5 ? valid_252 : _GEN_4628; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5666 = _T_5 ? valid_253 : _GEN_4629; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5667 = _T_5 ? valid_254 : _GEN_4630; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_5668 = _T_5 ? valid_255 : _GEN_4631; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire [19:0] _GEN_5669 = _T_5 ? tag_0 : _GEN_4632; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5670 = _T_5 ? tag_1 : _GEN_4633; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5671 = _T_5 ? tag_2 : _GEN_4634; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5672 = _T_5 ? tag_3 : _GEN_4635; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5673 = _T_5 ? tag_4 : _GEN_4636; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5674 = _T_5 ? tag_5 : _GEN_4637; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5675 = _T_5 ? tag_6 : _GEN_4638; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5676 = _T_5 ? tag_7 : _GEN_4639; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5677 = _T_5 ? tag_8 : _GEN_4640; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5678 = _T_5 ? tag_9 : _GEN_4641; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5679 = _T_5 ? tag_10 : _GEN_4642; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5680 = _T_5 ? tag_11 : _GEN_4643; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5681 = _T_5 ? tag_12 : _GEN_4644; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5682 = _T_5 ? tag_13 : _GEN_4645; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5683 = _T_5 ? tag_14 : _GEN_4646; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5684 = _T_5 ? tag_15 : _GEN_4647; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5685 = _T_5 ? tag_16 : _GEN_4648; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5686 = _T_5 ? tag_17 : _GEN_4649; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5687 = _T_5 ? tag_18 : _GEN_4650; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5688 = _T_5 ? tag_19 : _GEN_4651; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5689 = _T_5 ? tag_20 : _GEN_4652; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5690 = _T_5 ? tag_21 : _GEN_4653; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5691 = _T_5 ? tag_22 : _GEN_4654; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5692 = _T_5 ? tag_23 : _GEN_4655; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5693 = _T_5 ? tag_24 : _GEN_4656; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5694 = _T_5 ? tag_25 : _GEN_4657; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5695 = _T_5 ? tag_26 : _GEN_4658; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5696 = _T_5 ? tag_27 : _GEN_4659; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5697 = _T_5 ? tag_28 : _GEN_4660; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5698 = _T_5 ? tag_29 : _GEN_4661; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5699 = _T_5 ? tag_30 : _GEN_4662; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5700 = _T_5 ? tag_31 : _GEN_4663; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5701 = _T_5 ? tag_32 : _GEN_4664; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5702 = _T_5 ? tag_33 : _GEN_4665; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5703 = _T_5 ? tag_34 : _GEN_4666; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5704 = _T_5 ? tag_35 : _GEN_4667; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5705 = _T_5 ? tag_36 : _GEN_4668; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5706 = _T_5 ? tag_37 : _GEN_4669; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5707 = _T_5 ? tag_38 : _GEN_4670; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5708 = _T_5 ? tag_39 : _GEN_4671; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5709 = _T_5 ? tag_40 : _GEN_4672; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5710 = _T_5 ? tag_41 : _GEN_4673; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5711 = _T_5 ? tag_42 : _GEN_4674; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5712 = _T_5 ? tag_43 : _GEN_4675; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5713 = _T_5 ? tag_44 : _GEN_4676; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5714 = _T_5 ? tag_45 : _GEN_4677; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5715 = _T_5 ? tag_46 : _GEN_4678; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5716 = _T_5 ? tag_47 : _GEN_4679; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5717 = _T_5 ? tag_48 : _GEN_4680; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5718 = _T_5 ? tag_49 : _GEN_4681; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5719 = _T_5 ? tag_50 : _GEN_4682; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5720 = _T_5 ? tag_51 : _GEN_4683; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5721 = _T_5 ? tag_52 : _GEN_4684; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5722 = _T_5 ? tag_53 : _GEN_4685; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5723 = _T_5 ? tag_54 : _GEN_4686; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5724 = _T_5 ? tag_55 : _GEN_4687; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5725 = _T_5 ? tag_56 : _GEN_4688; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5726 = _T_5 ? tag_57 : _GEN_4689; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5727 = _T_5 ? tag_58 : _GEN_4690; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5728 = _T_5 ? tag_59 : _GEN_4691; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5729 = _T_5 ? tag_60 : _GEN_4692; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5730 = _T_5 ? tag_61 : _GEN_4693; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5731 = _T_5 ? tag_62 : _GEN_4694; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5732 = _T_5 ? tag_63 : _GEN_4695; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5733 = _T_5 ? tag_64 : _GEN_4696; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5734 = _T_5 ? tag_65 : _GEN_4697; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5735 = _T_5 ? tag_66 : _GEN_4698; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5736 = _T_5 ? tag_67 : _GEN_4699; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5737 = _T_5 ? tag_68 : _GEN_4700; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5738 = _T_5 ? tag_69 : _GEN_4701; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5739 = _T_5 ? tag_70 : _GEN_4702; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5740 = _T_5 ? tag_71 : _GEN_4703; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5741 = _T_5 ? tag_72 : _GEN_4704; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5742 = _T_5 ? tag_73 : _GEN_4705; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5743 = _T_5 ? tag_74 : _GEN_4706; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5744 = _T_5 ? tag_75 : _GEN_4707; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5745 = _T_5 ? tag_76 : _GEN_4708; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5746 = _T_5 ? tag_77 : _GEN_4709; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5747 = _T_5 ? tag_78 : _GEN_4710; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5748 = _T_5 ? tag_79 : _GEN_4711; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5749 = _T_5 ? tag_80 : _GEN_4712; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5750 = _T_5 ? tag_81 : _GEN_4713; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5751 = _T_5 ? tag_82 : _GEN_4714; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5752 = _T_5 ? tag_83 : _GEN_4715; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5753 = _T_5 ? tag_84 : _GEN_4716; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5754 = _T_5 ? tag_85 : _GEN_4717; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5755 = _T_5 ? tag_86 : _GEN_4718; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5756 = _T_5 ? tag_87 : _GEN_4719; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5757 = _T_5 ? tag_88 : _GEN_4720; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5758 = _T_5 ? tag_89 : _GEN_4721; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5759 = _T_5 ? tag_90 : _GEN_4722; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5760 = _T_5 ? tag_91 : _GEN_4723; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5761 = _T_5 ? tag_92 : _GEN_4724; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5762 = _T_5 ? tag_93 : _GEN_4725; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5763 = _T_5 ? tag_94 : _GEN_4726; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5764 = _T_5 ? tag_95 : _GEN_4727; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5765 = _T_5 ? tag_96 : _GEN_4728; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5766 = _T_5 ? tag_97 : _GEN_4729; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5767 = _T_5 ? tag_98 : _GEN_4730; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5768 = _T_5 ? tag_99 : _GEN_4731; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5769 = _T_5 ? tag_100 : _GEN_4732; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5770 = _T_5 ? tag_101 : _GEN_4733; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5771 = _T_5 ? tag_102 : _GEN_4734; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5772 = _T_5 ? tag_103 : _GEN_4735; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5773 = _T_5 ? tag_104 : _GEN_4736; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5774 = _T_5 ? tag_105 : _GEN_4737; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5775 = _T_5 ? tag_106 : _GEN_4738; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5776 = _T_5 ? tag_107 : _GEN_4739; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5777 = _T_5 ? tag_108 : _GEN_4740; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5778 = _T_5 ? tag_109 : _GEN_4741; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5779 = _T_5 ? tag_110 : _GEN_4742; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5780 = _T_5 ? tag_111 : _GEN_4743; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5781 = _T_5 ? tag_112 : _GEN_4744; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5782 = _T_5 ? tag_113 : _GEN_4745; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5783 = _T_5 ? tag_114 : _GEN_4746; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5784 = _T_5 ? tag_115 : _GEN_4747; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5785 = _T_5 ? tag_116 : _GEN_4748; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5786 = _T_5 ? tag_117 : _GEN_4749; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5787 = _T_5 ? tag_118 : _GEN_4750; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5788 = _T_5 ? tag_119 : _GEN_4751; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5789 = _T_5 ? tag_120 : _GEN_4752; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5790 = _T_5 ? tag_121 : _GEN_4753; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5791 = _T_5 ? tag_122 : _GEN_4754; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5792 = _T_5 ? tag_123 : _GEN_4755; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5793 = _T_5 ? tag_124 : _GEN_4756; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5794 = _T_5 ? tag_125 : _GEN_4757; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5795 = _T_5 ? tag_126 : _GEN_4758; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5796 = _T_5 ? tag_127 : _GEN_4759; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5797 = _T_5 ? tag_128 : _GEN_4760; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5798 = _T_5 ? tag_129 : _GEN_4761; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5799 = _T_5 ? tag_130 : _GEN_4762; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5800 = _T_5 ? tag_131 : _GEN_4763; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5801 = _T_5 ? tag_132 : _GEN_4764; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5802 = _T_5 ? tag_133 : _GEN_4765; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5803 = _T_5 ? tag_134 : _GEN_4766; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5804 = _T_5 ? tag_135 : _GEN_4767; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5805 = _T_5 ? tag_136 : _GEN_4768; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5806 = _T_5 ? tag_137 : _GEN_4769; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5807 = _T_5 ? tag_138 : _GEN_4770; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5808 = _T_5 ? tag_139 : _GEN_4771; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5809 = _T_5 ? tag_140 : _GEN_4772; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5810 = _T_5 ? tag_141 : _GEN_4773; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5811 = _T_5 ? tag_142 : _GEN_4774; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5812 = _T_5 ? tag_143 : _GEN_4775; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5813 = _T_5 ? tag_144 : _GEN_4776; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5814 = _T_5 ? tag_145 : _GEN_4777; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5815 = _T_5 ? tag_146 : _GEN_4778; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5816 = _T_5 ? tag_147 : _GEN_4779; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5817 = _T_5 ? tag_148 : _GEN_4780; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5818 = _T_5 ? tag_149 : _GEN_4781; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5819 = _T_5 ? tag_150 : _GEN_4782; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5820 = _T_5 ? tag_151 : _GEN_4783; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5821 = _T_5 ? tag_152 : _GEN_4784; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5822 = _T_5 ? tag_153 : _GEN_4785; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5823 = _T_5 ? tag_154 : _GEN_4786; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5824 = _T_5 ? tag_155 : _GEN_4787; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5825 = _T_5 ? tag_156 : _GEN_4788; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5826 = _T_5 ? tag_157 : _GEN_4789; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5827 = _T_5 ? tag_158 : _GEN_4790; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5828 = _T_5 ? tag_159 : _GEN_4791; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5829 = _T_5 ? tag_160 : _GEN_4792; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5830 = _T_5 ? tag_161 : _GEN_4793; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5831 = _T_5 ? tag_162 : _GEN_4794; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5832 = _T_5 ? tag_163 : _GEN_4795; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5833 = _T_5 ? tag_164 : _GEN_4796; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5834 = _T_5 ? tag_165 : _GEN_4797; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5835 = _T_5 ? tag_166 : _GEN_4798; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5836 = _T_5 ? tag_167 : _GEN_4799; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5837 = _T_5 ? tag_168 : _GEN_4800; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5838 = _T_5 ? tag_169 : _GEN_4801; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5839 = _T_5 ? tag_170 : _GEN_4802; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5840 = _T_5 ? tag_171 : _GEN_4803; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5841 = _T_5 ? tag_172 : _GEN_4804; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5842 = _T_5 ? tag_173 : _GEN_4805; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5843 = _T_5 ? tag_174 : _GEN_4806; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5844 = _T_5 ? tag_175 : _GEN_4807; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5845 = _T_5 ? tag_176 : _GEN_4808; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5846 = _T_5 ? tag_177 : _GEN_4809; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5847 = _T_5 ? tag_178 : _GEN_4810; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5848 = _T_5 ? tag_179 : _GEN_4811; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5849 = _T_5 ? tag_180 : _GEN_4812; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5850 = _T_5 ? tag_181 : _GEN_4813; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5851 = _T_5 ? tag_182 : _GEN_4814; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5852 = _T_5 ? tag_183 : _GEN_4815; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5853 = _T_5 ? tag_184 : _GEN_4816; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5854 = _T_5 ? tag_185 : _GEN_4817; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5855 = _T_5 ? tag_186 : _GEN_4818; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5856 = _T_5 ? tag_187 : _GEN_4819; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5857 = _T_5 ? tag_188 : _GEN_4820; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5858 = _T_5 ? tag_189 : _GEN_4821; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5859 = _T_5 ? tag_190 : _GEN_4822; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5860 = _T_5 ? tag_191 : _GEN_4823; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5861 = _T_5 ? tag_192 : _GEN_4824; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5862 = _T_5 ? tag_193 : _GEN_4825; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5863 = _T_5 ? tag_194 : _GEN_4826; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5864 = _T_5 ? tag_195 : _GEN_4827; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5865 = _T_5 ? tag_196 : _GEN_4828; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5866 = _T_5 ? tag_197 : _GEN_4829; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5867 = _T_5 ? tag_198 : _GEN_4830; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5868 = _T_5 ? tag_199 : _GEN_4831; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5869 = _T_5 ? tag_200 : _GEN_4832; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5870 = _T_5 ? tag_201 : _GEN_4833; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5871 = _T_5 ? tag_202 : _GEN_4834; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5872 = _T_5 ? tag_203 : _GEN_4835; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5873 = _T_5 ? tag_204 : _GEN_4836; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5874 = _T_5 ? tag_205 : _GEN_4837; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5875 = _T_5 ? tag_206 : _GEN_4838; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5876 = _T_5 ? tag_207 : _GEN_4839; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5877 = _T_5 ? tag_208 : _GEN_4840; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5878 = _T_5 ? tag_209 : _GEN_4841; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5879 = _T_5 ? tag_210 : _GEN_4842; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5880 = _T_5 ? tag_211 : _GEN_4843; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5881 = _T_5 ? tag_212 : _GEN_4844; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5882 = _T_5 ? tag_213 : _GEN_4845; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5883 = _T_5 ? tag_214 : _GEN_4846; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5884 = _T_5 ? tag_215 : _GEN_4847; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5885 = _T_5 ? tag_216 : _GEN_4848; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5886 = _T_5 ? tag_217 : _GEN_4849; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5887 = _T_5 ? tag_218 : _GEN_4850; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5888 = _T_5 ? tag_219 : _GEN_4851; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5889 = _T_5 ? tag_220 : _GEN_4852; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5890 = _T_5 ? tag_221 : _GEN_4853; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5891 = _T_5 ? tag_222 : _GEN_4854; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5892 = _T_5 ? tag_223 : _GEN_4855; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5893 = _T_5 ? tag_224 : _GEN_4856; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5894 = _T_5 ? tag_225 : _GEN_4857; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5895 = _T_5 ? tag_226 : _GEN_4858; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5896 = _T_5 ? tag_227 : _GEN_4859; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5897 = _T_5 ? tag_228 : _GEN_4860; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5898 = _T_5 ? tag_229 : _GEN_4861; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5899 = _T_5 ? tag_230 : _GEN_4862; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5900 = _T_5 ? tag_231 : _GEN_4863; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5901 = _T_5 ? tag_232 : _GEN_4864; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5902 = _T_5 ? tag_233 : _GEN_4865; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5903 = _T_5 ? tag_234 : _GEN_4866; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5904 = _T_5 ? tag_235 : _GEN_4867; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5905 = _T_5 ? tag_236 : _GEN_4868; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5906 = _T_5 ? tag_237 : _GEN_4869; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5907 = _T_5 ? tag_238 : _GEN_4870; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5908 = _T_5 ? tag_239 : _GEN_4871; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5909 = _T_5 ? tag_240 : _GEN_4872; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5910 = _T_5 ? tag_241 : _GEN_4873; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5911 = _T_5 ? tag_242 : _GEN_4874; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5912 = _T_5 ? tag_243 : _GEN_4875; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5913 = _T_5 ? tag_244 : _GEN_4876; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5914 = _T_5 ? tag_245 : _GEN_4877; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5915 = _T_5 ? tag_246 : _GEN_4878; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5916 = _T_5 ? tag_247 : _GEN_4879; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5917 = _T_5 ? tag_248 : _GEN_4880; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5918 = _T_5 ? tag_249 : _GEN_4881; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5919 = _T_5 ? tag_250 : _GEN_4882; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5920 = _T_5 ? tag_251 : _GEN_4883; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5921 = _T_5 ? tag_252 : _GEN_4884; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5922 = _T_5 ? tag_253 : _GEN_4885; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5923 = _T_5 ? tag_254 : _GEN_4886; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_5924 = _T_5 ? tag_255 : _GEN_4887; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire  _GEN_5925 = _T_5 ? dirty_0 : _GEN_4888; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5926 = _T_5 ? dirty_1 : _GEN_4889; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5927 = _T_5 ? dirty_2 : _GEN_4890; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5928 = _T_5 ? dirty_3 : _GEN_4891; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5929 = _T_5 ? dirty_4 : _GEN_4892; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5930 = _T_5 ? dirty_5 : _GEN_4893; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5931 = _T_5 ? dirty_6 : _GEN_4894; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5932 = _T_5 ? dirty_7 : _GEN_4895; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5933 = _T_5 ? dirty_8 : _GEN_4896; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5934 = _T_5 ? dirty_9 : _GEN_4897; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5935 = _T_5 ? dirty_10 : _GEN_4898; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5936 = _T_5 ? dirty_11 : _GEN_4899; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5937 = _T_5 ? dirty_12 : _GEN_4900; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5938 = _T_5 ? dirty_13 : _GEN_4901; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5939 = _T_5 ? dirty_14 : _GEN_4902; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5940 = _T_5 ? dirty_15 : _GEN_4903; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5941 = _T_5 ? dirty_16 : _GEN_4904; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5942 = _T_5 ? dirty_17 : _GEN_4905; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5943 = _T_5 ? dirty_18 : _GEN_4906; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5944 = _T_5 ? dirty_19 : _GEN_4907; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5945 = _T_5 ? dirty_20 : _GEN_4908; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5946 = _T_5 ? dirty_21 : _GEN_4909; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5947 = _T_5 ? dirty_22 : _GEN_4910; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5948 = _T_5 ? dirty_23 : _GEN_4911; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5949 = _T_5 ? dirty_24 : _GEN_4912; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5950 = _T_5 ? dirty_25 : _GEN_4913; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5951 = _T_5 ? dirty_26 : _GEN_4914; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5952 = _T_5 ? dirty_27 : _GEN_4915; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5953 = _T_5 ? dirty_28 : _GEN_4916; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5954 = _T_5 ? dirty_29 : _GEN_4917; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5955 = _T_5 ? dirty_30 : _GEN_4918; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5956 = _T_5 ? dirty_31 : _GEN_4919; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5957 = _T_5 ? dirty_32 : _GEN_4920; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5958 = _T_5 ? dirty_33 : _GEN_4921; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5959 = _T_5 ? dirty_34 : _GEN_4922; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5960 = _T_5 ? dirty_35 : _GEN_4923; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5961 = _T_5 ? dirty_36 : _GEN_4924; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5962 = _T_5 ? dirty_37 : _GEN_4925; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5963 = _T_5 ? dirty_38 : _GEN_4926; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5964 = _T_5 ? dirty_39 : _GEN_4927; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5965 = _T_5 ? dirty_40 : _GEN_4928; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5966 = _T_5 ? dirty_41 : _GEN_4929; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5967 = _T_5 ? dirty_42 : _GEN_4930; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5968 = _T_5 ? dirty_43 : _GEN_4931; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5969 = _T_5 ? dirty_44 : _GEN_4932; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5970 = _T_5 ? dirty_45 : _GEN_4933; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5971 = _T_5 ? dirty_46 : _GEN_4934; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5972 = _T_5 ? dirty_47 : _GEN_4935; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5973 = _T_5 ? dirty_48 : _GEN_4936; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5974 = _T_5 ? dirty_49 : _GEN_4937; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5975 = _T_5 ? dirty_50 : _GEN_4938; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5976 = _T_5 ? dirty_51 : _GEN_4939; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5977 = _T_5 ? dirty_52 : _GEN_4940; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5978 = _T_5 ? dirty_53 : _GEN_4941; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5979 = _T_5 ? dirty_54 : _GEN_4942; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5980 = _T_5 ? dirty_55 : _GEN_4943; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5981 = _T_5 ? dirty_56 : _GEN_4944; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5982 = _T_5 ? dirty_57 : _GEN_4945; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5983 = _T_5 ? dirty_58 : _GEN_4946; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5984 = _T_5 ? dirty_59 : _GEN_4947; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5985 = _T_5 ? dirty_60 : _GEN_4948; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5986 = _T_5 ? dirty_61 : _GEN_4949; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5987 = _T_5 ? dirty_62 : _GEN_4950; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5988 = _T_5 ? dirty_63 : _GEN_4951; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5989 = _T_5 ? dirty_64 : _GEN_4952; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5990 = _T_5 ? dirty_65 : _GEN_4953; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5991 = _T_5 ? dirty_66 : _GEN_4954; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5992 = _T_5 ? dirty_67 : _GEN_4955; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5993 = _T_5 ? dirty_68 : _GEN_4956; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5994 = _T_5 ? dirty_69 : _GEN_4957; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5995 = _T_5 ? dirty_70 : _GEN_4958; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5996 = _T_5 ? dirty_71 : _GEN_4959; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5997 = _T_5 ? dirty_72 : _GEN_4960; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5998 = _T_5 ? dirty_73 : _GEN_4961; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_5999 = _T_5 ? dirty_74 : _GEN_4962; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6000 = _T_5 ? dirty_75 : _GEN_4963; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6001 = _T_5 ? dirty_76 : _GEN_4964; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6002 = _T_5 ? dirty_77 : _GEN_4965; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6003 = _T_5 ? dirty_78 : _GEN_4966; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6004 = _T_5 ? dirty_79 : _GEN_4967; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6005 = _T_5 ? dirty_80 : _GEN_4968; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6006 = _T_5 ? dirty_81 : _GEN_4969; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6007 = _T_5 ? dirty_82 : _GEN_4970; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6008 = _T_5 ? dirty_83 : _GEN_4971; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6009 = _T_5 ? dirty_84 : _GEN_4972; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6010 = _T_5 ? dirty_85 : _GEN_4973; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6011 = _T_5 ? dirty_86 : _GEN_4974; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6012 = _T_5 ? dirty_87 : _GEN_4975; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6013 = _T_5 ? dirty_88 : _GEN_4976; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6014 = _T_5 ? dirty_89 : _GEN_4977; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6015 = _T_5 ? dirty_90 : _GEN_4978; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6016 = _T_5 ? dirty_91 : _GEN_4979; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6017 = _T_5 ? dirty_92 : _GEN_4980; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6018 = _T_5 ? dirty_93 : _GEN_4981; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6019 = _T_5 ? dirty_94 : _GEN_4982; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6020 = _T_5 ? dirty_95 : _GEN_4983; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6021 = _T_5 ? dirty_96 : _GEN_4984; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6022 = _T_5 ? dirty_97 : _GEN_4985; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6023 = _T_5 ? dirty_98 : _GEN_4986; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6024 = _T_5 ? dirty_99 : _GEN_4987; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6025 = _T_5 ? dirty_100 : _GEN_4988; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6026 = _T_5 ? dirty_101 : _GEN_4989; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6027 = _T_5 ? dirty_102 : _GEN_4990; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6028 = _T_5 ? dirty_103 : _GEN_4991; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6029 = _T_5 ? dirty_104 : _GEN_4992; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6030 = _T_5 ? dirty_105 : _GEN_4993; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6031 = _T_5 ? dirty_106 : _GEN_4994; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6032 = _T_5 ? dirty_107 : _GEN_4995; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6033 = _T_5 ? dirty_108 : _GEN_4996; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6034 = _T_5 ? dirty_109 : _GEN_4997; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6035 = _T_5 ? dirty_110 : _GEN_4998; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6036 = _T_5 ? dirty_111 : _GEN_4999; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6037 = _T_5 ? dirty_112 : _GEN_5000; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6038 = _T_5 ? dirty_113 : _GEN_5001; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6039 = _T_5 ? dirty_114 : _GEN_5002; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6040 = _T_5 ? dirty_115 : _GEN_5003; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6041 = _T_5 ? dirty_116 : _GEN_5004; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6042 = _T_5 ? dirty_117 : _GEN_5005; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6043 = _T_5 ? dirty_118 : _GEN_5006; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6044 = _T_5 ? dirty_119 : _GEN_5007; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6045 = _T_5 ? dirty_120 : _GEN_5008; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6046 = _T_5 ? dirty_121 : _GEN_5009; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6047 = _T_5 ? dirty_122 : _GEN_5010; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6048 = _T_5 ? dirty_123 : _GEN_5011; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6049 = _T_5 ? dirty_124 : _GEN_5012; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6050 = _T_5 ? dirty_125 : _GEN_5013; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6051 = _T_5 ? dirty_126 : _GEN_5014; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6052 = _T_5 ? dirty_127 : _GEN_5015; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6053 = _T_5 ? dirty_128 : _GEN_5016; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6054 = _T_5 ? dirty_129 : _GEN_5017; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6055 = _T_5 ? dirty_130 : _GEN_5018; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6056 = _T_5 ? dirty_131 : _GEN_5019; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6057 = _T_5 ? dirty_132 : _GEN_5020; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6058 = _T_5 ? dirty_133 : _GEN_5021; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6059 = _T_5 ? dirty_134 : _GEN_5022; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6060 = _T_5 ? dirty_135 : _GEN_5023; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6061 = _T_5 ? dirty_136 : _GEN_5024; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6062 = _T_5 ? dirty_137 : _GEN_5025; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6063 = _T_5 ? dirty_138 : _GEN_5026; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6064 = _T_5 ? dirty_139 : _GEN_5027; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6065 = _T_5 ? dirty_140 : _GEN_5028; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6066 = _T_5 ? dirty_141 : _GEN_5029; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6067 = _T_5 ? dirty_142 : _GEN_5030; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6068 = _T_5 ? dirty_143 : _GEN_5031; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6069 = _T_5 ? dirty_144 : _GEN_5032; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6070 = _T_5 ? dirty_145 : _GEN_5033; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6071 = _T_5 ? dirty_146 : _GEN_5034; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6072 = _T_5 ? dirty_147 : _GEN_5035; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6073 = _T_5 ? dirty_148 : _GEN_5036; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6074 = _T_5 ? dirty_149 : _GEN_5037; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6075 = _T_5 ? dirty_150 : _GEN_5038; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6076 = _T_5 ? dirty_151 : _GEN_5039; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6077 = _T_5 ? dirty_152 : _GEN_5040; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6078 = _T_5 ? dirty_153 : _GEN_5041; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6079 = _T_5 ? dirty_154 : _GEN_5042; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6080 = _T_5 ? dirty_155 : _GEN_5043; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6081 = _T_5 ? dirty_156 : _GEN_5044; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6082 = _T_5 ? dirty_157 : _GEN_5045; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6083 = _T_5 ? dirty_158 : _GEN_5046; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6084 = _T_5 ? dirty_159 : _GEN_5047; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6085 = _T_5 ? dirty_160 : _GEN_5048; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6086 = _T_5 ? dirty_161 : _GEN_5049; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6087 = _T_5 ? dirty_162 : _GEN_5050; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6088 = _T_5 ? dirty_163 : _GEN_5051; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6089 = _T_5 ? dirty_164 : _GEN_5052; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6090 = _T_5 ? dirty_165 : _GEN_5053; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6091 = _T_5 ? dirty_166 : _GEN_5054; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6092 = _T_5 ? dirty_167 : _GEN_5055; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6093 = _T_5 ? dirty_168 : _GEN_5056; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6094 = _T_5 ? dirty_169 : _GEN_5057; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6095 = _T_5 ? dirty_170 : _GEN_5058; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6096 = _T_5 ? dirty_171 : _GEN_5059; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6097 = _T_5 ? dirty_172 : _GEN_5060; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6098 = _T_5 ? dirty_173 : _GEN_5061; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6099 = _T_5 ? dirty_174 : _GEN_5062; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6100 = _T_5 ? dirty_175 : _GEN_5063; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6101 = _T_5 ? dirty_176 : _GEN_5064; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6102 = _T_5 ? dirty_177 : _GEN_5065; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6103 = _T_5 ? dirty_178 : _GEN_5066; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6104 = _T_5 ? dirty_179 : _GEN_5067; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6105 = _T_5 ? dirty_180 : _GEN_5068; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6106 = _T_5 ? dirty_181 : _GEN_5069; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6107 = _T_5 ? dirty_182 : _GEN_5070; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6108 = _T_5 ? dirty_183 : _GEN_5071; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6109 = _T_5 ? dirty_184 : _GEN_5072; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6110 = _T_5 ? dirty_185 : _GEN_5073; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6111 = _T_5 ? dirty_186 : _GEN_5074; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6112 = _T_5 ? dirty_187 : _GEN_5075; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6113 = _T_5 ? dirty_188 : _GEN_5076; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6114 = _T_5 ? dirty_189 : _GEN_5077; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6115 = _T_5 ? dirty_190 : _GEN_5078; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6116 = _T_5 ? dirty_191 : _GEN_5079; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6117 = _T_5 ? dirty_192 : _GEN_5080; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6118 = _T_5 ? dirty_193 : _GEN_5081; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6119 = _T_5 ? dirty_194 : _GEN_5082; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6120 = _T_5 ? dirty_195 : _GEN_5083; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6121 = _T_5 ? dirty_196 : _GEN_5084; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6122 = _T_5 ? dirty_197 : _GEN_5085; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6123 = _T_5 ? dirty_198 : _GEN_5086; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6124 = _T_5 ? dirty_199 : _GEN_5087; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6125 = _T_5 ? dirty_200 : _GEN_5088; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6126 = _T_5 ? dirty_201 : _GEN_5089; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6127 = _T_5 ? dirty_202 : _GEN_5090; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6128 = _T_5 ? dirty_203 : _GEN_5091; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6129 = _T_5 ? dirty_204 : _GEN_5092; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6130 = _T_5 ? dirty_205 : _GEN_5093; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6131 = _T_5 ? dirty_206 : _GEN_5094; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6132 = _T_5 ? dirty_207 : _GEN_5095; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6133 = _T_5 ? dirty_208 : _GEN_5096; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6134 = _T_5 ? dirty_209 : _GEN_5097; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6135 = _T_5 ? dirty_210 : _GEN_5098; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6136 = _T_5 ? dirty_211 : _GEN_5099; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6137 = _T_5 ? dirty_212 : _GEN_5100; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6138 = _T_5 ? dirty_213 : _GEN_5101; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6139 = _T_5 ? dirty_214 : _GEN_5102; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6140 = _T_5 ? dirty_215 : _GEN_5103; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6141 = _T_5 ? dirty_216 : _GEN_5104; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6142 = _T_5 ? dirty_217 : _GEN_5105; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6143 = _T_5 ? dirty_218 : _GEN_5106; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6144 = _T_5 ? dirty_219 : _GEN_5107; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6145 = _T_5 ? dirty_220 : _GEN_5108; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6146 = _T_5 ? dirty_221 : _GEN_5109; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6147 = _T_5 ? dirty_222 : _GEN_5110; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6148 = _T_5 ? dirty_223 : _GEN_5111; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6149 = _T_5 ? dirty_224 : _GEN_5112; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6150 = _T_5 ? dirty_225 : _GEN_5113; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6151 = _T_5 ? dirty_226 : _GEN_5114; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6152 = _T_5 ? dirty_227 : _GEN_5115; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6153 = _T_5 ? dirty_228 : _GEN_5116; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6154 = _T_5 ? dirty_229 : _GEN_5117; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6155 = _T_5 ? dirty_230 : _GEN_5118; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6156 = _T_5 ? dirty_231 : _GEN_5119; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6157 = _T_5 ? dirty_232 : _GEN_5120; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6158 = _T_5 ? dirty_233 : _GEN_5121; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6159 = _T_5 ? dirty_234 : _GEN_5122; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6160 = _T_5 ? dirty_235 : _GEN_5123; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6161 = _T_5 ? dirty_236 : _GEN_5124; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6162 = _T_5 ? dirty_237 : _GEN_5125; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6163 = _T_5 ? dirty_238 : _GEN_5126; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6164 = _T_5 ? dirty_239 : _GEN_5127; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6165 = _T_5 ? dirty_240 : _GEN_5128; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6166 = _T_5 ? dirty_241 : _GEN_5129; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6167 = _T_5 ? dirty_242 : _GEN_5130; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6168 = _T_5 ? dirty_243 : _GEN_5131; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6169 = _T_5 ? dirty_244 : _GEN_5132; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6170 = _T_5 ? dirty_245 : _GEN_5133; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6171 = _T_5 ? dirty_246 : _GEN_5134; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6172 = _T_5 ? dirty_247 : _GEN_5135; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6173 = _T_5 ? dirty_248 : _GEN_5136; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6174 = _T_5 ? dirty_249 : _GEN_5137; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6175 = _T_5 ? dirty_250 : _GEN_5138; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6176 = _T_5 ? dirty_251 : _GEN_5139; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6177 = _T_5 ? dirty_252 : _GEN_5140; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6178 = _T_5 ? dirty_253 : _GEN_5141; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6179 = _T_5 ? dirty_254 : _GEN_5142; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6180 = _T_5 ? dirty_255 : _GEN_5143; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire [3:0] _GEN_6181 = _T_5 ? offset_0 : _GEN_5144; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6182 = _T_5 ? offset_1 : _GEN_5145; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6183 = _T_5 ? offset_2 : _GEN_5146; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6184 = _T_5 ? offset_3 : _GEN_5147; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6185 = _T_5 ? offset_4 : _GEN_5148; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6186 = _T_5 ? offset_5 : _GEN_5149; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6187 = _T_5 ? offset_6 : _GEN_5150; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6188 = _T_5 ? offset_7 : _GEN_5151; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6189 = _T_5 ? offset_8 : _GEN_5152; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6190 = _T_5 ? offset_9 : _GEN_5153; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6191 = _T_5 ? offset_10 : _GEN_5154; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6192 = _T_5 ? offset_11 : _GEN_5155; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6193 = _T_5 ? offset_12 : _GEN_5156; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6194 = _T_5 ? offset_13 : _GEN_5157; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6195 = _T_5 ? offset_14 : _GEN_5158; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6196 = _T_5 ? offset_15 : _GEN_5159; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6197 = _T_5 ? offset_16 : _GEN_5160; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6198 = _T_5 ? offset_17 : _GEN_5161; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6199 = _T_5 ? offset_18 : _GEN_5162; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6200 = _T_5 ? offset_19 : _GEN_5163; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6201 = _T_5 ? offset_20 : _GEN_5164; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6202 = _T_5 ? offset_21 : _GEN_5165; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6203 = _T_5 ? offset_22 : _GEN_5166; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6204 = _T_5 ? offset_23 : _GEN_5167; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6205 = _T_5 ? offset_24 : _GEN_5168; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6206 = _T_5 ? offset_25 : _GEN_5169; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6207 = _T_5 ? offset_26 : _GEN_5170; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6208 = _T_5 ? offset_27 : _GEN_5171; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6209 = _T_5 ? offset_28 : _GEN_5172; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6210 = _T_5 ? offset_29 : _GEN_5173; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6211 = _T_5 ? offset_30 : _GEN_5174; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6212 = _T_5 ? offset_31 : _GEN_5175; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6213 = _T_5 ? offset_32 : _GEN_5176; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6214 = _T_5 ? offset_33 : _GEN_5177; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6215 = _T_5 ? offset_34 : _GEN_5178; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6216 = _T_5 ? offset_35 : _GEN_5179; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6217 = _T_5 ? offset_36 : _GEN_5180; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6218 = _T_5 ? offset_37 : _GEN_5181; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6219 = _T_5 ? offset_38 : _GEN_5182; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6220 = _T_5 ? offset_39 : _GEN_5183; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6221 = _T_5 ? offset_40 : _GEN_5184; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6222 = _T_5 ? offset_41 : _GEN_5185; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6223 = _T_5 ? offset_42 : _GEN_5186; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6224 = _T_5 ? offset_43 : _GEN_5187; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6225 = _T_5 ? offset_44 : _GEN_5188; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6226 = _T_5 ? offset_45 : _GEN_5189; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6227 = _T_5 ? offset_46 : _GEN_5190; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6228 = _T_5 ? offset_47 : _GEN_5191; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6229 = _T_5 ? offset_48 : _GEN_5192; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6230 = _T_5 ? offset_49 : _GEN_5193; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6231 = _T_5 ? offset_50 : _GEN_5194; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6232 = _T_5 ? offset_51 : _GEN_5195; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6233 = _T_5 ? offset_52 : _GEN_5196; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6234 = _T_5 ? offset_53 : _GEN_5197; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6235 = _T_5 ? offset_54 : _GEN_5198; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6236 = _T_5 ? offset_55 : _GEN_5199; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6237 = _T_5 ? offset_56 : _GEN_5200; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6238 = _T_5 ? offset_57 : _GEN_5201; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6239 = _T_5 ? offset_58 : _GEN_5202; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6240 = _T_5 ? offset_59 : _GEN_5203; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6241 = _T_5 ? offset_60 : _GEN_5204; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6242 = _T_5 ? offset_61 : _GEN_5205; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6243 = _T_5 ? offset_62 : _GEN_5206; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6244 = _T_5 ? offset_63 : _GEN_5207; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6245 = _T_5 ? offset_64 : _GEN_5208; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6246 = _T_5 ? offset_65 : _GEN_5209; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6247 = _T_5 ? offset_66 : _GEN_5210; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6248 = _T_5 ? offset_67 : _GEN_5211; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6249 = _T_5 ? offset_68 : _GEN_5212; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6250 = _T_5 ? offset_69 : _GEN_5213; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6251 = _T_5 ? offset_70 : _GEN_5214; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6252 = _T_5 ? offset_71 : _GEN_5215; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6253 = _T_5 ? offset_72 : _GEN_5216; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6254 = _T_5 ? offset_73 : _GEN_5217; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6255 = _T_5 ? offset_74 : _GEN_5218; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6256 = _T_5 ? offset_75 : _GEN_5219; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6257 = _T_5 ? offset_76 : _GEN_5220; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6258 = _T_5 ? offset_77 : _GEN_5221; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6259 = _T_5 ? offset_78 : _GEN_5222; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6260 = _T_5 ? offset_79 : _GEN_5223; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6261 = _T_5 ? offset_80 : _GEN_5224; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6262 = _T_5 ? offset_81 : _GEN_5225; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6263 = _T_5 ? offset_82 : _GEN_5226; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6264 = _T_5 ? offset_83 : _GEN_5227; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6265 = _T_5 ? offset_84 : _GEN_5228; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6266 = _T_5 ? offset_85 : _GEN_5229; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6267 = _T_5 ? offset_86 : _GEN_5230; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6268 = _T_5 ? offset_87 : _GEN_5231; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6269 = _T_5 ? offset_88 : _GEN_5232; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6270 = _T_5 ? offset_89 : _GEN_5233; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6271 = _T_5 ? offset_90 : _GEN_5234; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6272 = _T_5 ? offset_91 : _GEN_5235; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6273 = _T_5 ? offset_92 : _GEN_5236; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6274 = _T_5 ? offset_93 : _GEN_5237; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6275 = _T_5 ? offset_94 : _GEN_5238; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6276 = _T_5 ? offset_95 : _GEN_5239; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6277 = _T_5 ? offset_96 : _GEN_5240; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6278 = _T_5 ? offset_97 : _GEN_5241; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6279 = _T_5 ? offset_98 : _GEN_5242; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6280 = _T_5 ? offset_99 : _GEN_5243; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6281 = _T_5 ? offset_100 : _GEN_5244; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6282 = _T_5 ? offset_101 : _GEN_5245; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6283 = _T_5 ? offset_102 : _GEN_5246; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6284 = _T_5 ? offset_103 : _GEN_5247; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6285 = _T_5 ? offset_104 : _GEN_5248; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6286 = _T_5 ? offset_105 : _GEN_5249; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6287 = _T_5 ? offset_106 : _GEN_5250; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6288 = _T_5 ? offset_107 : _GEN_5251; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6289 = _T_5 ? offset_108 : _GEN_5252; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6290 = _T_5 ? offset_109 : _GEN_5253; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6291 = _T_5 ? offset_110 : _GEN_5254; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6292 = _T_5 ? offset_111 : _GEN_5255; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6293 = _T_5 ? offset_112 : _GEN_5256; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6294 = _T_5 ? offset_113 : _GEN_5257; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6295 = _T_5 ? offset_114 : _GEN_5258; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6296 = _T_5 ? offset_115 : _GEN_5259; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6297 = _T_5 ? offset_116 : _GEN_5260; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6298 = _T_5 ? offset_117 : _GEN_5261; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6299 = _T_5 ? offset_118 : _GEN_5262; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6300 = _T_5 ? offset_119 : _GEN_5263; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6301 = _T_5 ? offset_120 : _GEN_5264; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6302 = _T_5 ? offset_121 : _GEN_5265; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6303 = _T_5 ? offset_122 : _GEN_5266; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6304 = _T_5 ? offset_123 : _GEN_5267; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6305 = _T_5 ? offset_124 : _GEN_5268; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6306 = _T_5 ? offset_125 : _GEN_5269; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6307 = _T_5 ? offset_126 : _GEN_5270; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6308 = _T_5 ? offset_127 : _GEN_5271; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6309 = _T_5 ? offset_128 : _GEN_5272; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6310 = _T_5 ? offset_129 : _GEN_5273; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6311 = _T_5 ? offset_130 : _GEN_5274; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6312 = _T_5 ? offset_131 : _GEN_5275; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6313 = _T_5 ? offset_132 : _GEN_5276; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6314 = _T_5 ? offset_133 : _GEN_5277; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6315 = _T_5 ? offset_134 : _GEN_5278; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6316 = _T_5 ? offset_135 : _GEN_5279; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6317 = _T_5 ? offset_136 : _GEN_5280; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6318 = _T_5 ? offset_137 : _GEN_5281; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6319 = _T_5 ? offset_138 : _GEN_5282; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6320 = _T_5 ? offset_139 : _GEN_5283; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6321 = _T_5 ? offset_140 : _GEN_5284; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6322 = _T_5 ? offset_141 : _GEN_5285; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6323 = _T_5 ? offset_142 : _GEN_5286; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6324 = _T_5 ? offset_143 : _GEN_5287; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6325 = _T_5 ? offset_144 : _GEN_5288; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6326 = _T_5 ? offset_145 : _GEN_5289; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6327 = _T_5 ? offset_146 : _GEN_5290; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6328 = _T_5 ? offset_147 : _GEN_5291; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6329 = _T_5 ? offset_148 : _GEN_5292; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6330 = _T_5 ? offset_149 : _GEN_5293; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6331 = _T_5 ? offset_150 : _GEN_5294; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6332 = _T_5 ? offset_151 : _GEN_5295; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6333 = _T_5 ? offset_152 : _GEN_5296; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6334 = _T_5 ? offset_153 : _GEN_5297; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6335 = _T_5 ? offset_154 : _GEN_5298; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6336 = _T_5 ? offset_155 : _GEN_5299; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6337 = _T_5 ? offset_156 : _GEN_5300; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6338 = _T_5 ? offset_157 : _GEN_5301; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6339 = _T_5 ? offset_158 : _GEN_5302; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6340 = _T_5 ? offset_159 : _GEN_5303; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6341 = _T_5 ? offset_160 : _GEN_5304; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6342 = _T_5 ? offset_161 : _GEN_5305; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6343 = _T_5 ? offset_162 : _GEN_5306; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6344 = _T_5 ? offset_163 : _GEN_5307; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6345 = _T_5 ? offset_164 : _GEN_5308; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6346 = _T_5 ? offset_165 : _GEN_5309; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6347 = _T_5 ? offset_166 : _GEN_5310; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6348 = _T_5 ? offset_167 : _GEN_5311; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6349 = _T_5 ? offset_168 : _GEN_5312; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6350 = _T_5 ? offset_169 : _GEN_5313; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6351 = _T_5 ? offset_170 : _GEN_5314; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6352 = _T_5 ? offset_171 : _GEN_5315; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6353 = _T_5 ? offset_172 : _GEN_5316; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6354 = _T_5 ? offset_173 : _GEN_5317; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6355 = _T_5 ? offset_174 : _GEN_5318; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6356 = _T_5 ? offset_175 : _GEN_5319; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6357 = _T_5 ? offset_176 : _GEN_5320; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6358 = _T_5 ? offset_177 : _GEN_5321; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6359 = _T_5 ? offset_178 : _GEN_5322; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6360 = _T_5 ? offset_179 : _GEN_5323; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6361 = _T_5 ? offset_180 : _GEN_5324; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6362 = _T_5 ? offset_181 : _GEN_5325; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6363 = _T_5 ? offset_182 : _GEN_5326; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6364 = _T_5 ? offset_183 : _GEN_5327; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6365 = _T_5 ? offset_184 : _GEN_5328; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6366 = _T_5 ? offset_185 : _GEN_5329; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6367 = _T_5 ? offset_186 : _GEN_5330; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6368 = _T_5 ? offset_187 : _GEN_5331; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6369 = _T_5 ? offset_188 : _GEN_5332; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6370 = _T_5 ? offset_189 : _GEN_5333; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6371 = _T_5 ? offset_190 : _GEN_5334; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6372 = _T_5 ? offset_191 : _GEN_5335; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6373 = _T_5 ? offset_192 : _GEN_5336; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6374 = _T_5 ? offset_193 : _GEN_5337; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6375 = _T_5 ? offset_194 : _GEN_5338; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6376 = _T_5 ? offset_195 : _GEN_5339; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6377 = _T_5 ? offset_196 : _GEN_5340; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6378 = _T_5 ? offset_197 : _GEN_5341; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6379 = _T_5 ? offset_198 : _GEN_5342; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6380 = _T_5 ? offset_199 : _GEN_5343; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6381 = _T_5 ? offset_200 : _GEN_5344; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6382 = _T_5 ? offset_201 : _GEN_5345; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6383 = _T_5 ? offset_202 : _GEN_5346; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6384 = _T_5 ? offset_203 : _GEN_5347; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6385 = _T_5 ? offset_204 : _GEN_5348; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6386 = _T_5 ? offset_205 : _GEN_5349; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6387 = _T_5 ? offset_206 : _GEN_5350; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6388 = _T_5 ? offset_207 : _GEN_5351; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6389 = _T_5 ? offset_208 : _GEN_5352; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6390 = _T_5 ? offset_209 : _GEN_5353; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6391 = _T_5 ? offset_210 : _GEN_5354; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6392 = _T_5 ? offset_211 : _GEN_5355; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6393 = _T_5 ? offset_212 : _GEN_5356; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6394 = _T_5 ? offset_213 : _GEN_5357; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6395 = _T_5 ? offset_214 : _GEN_5358; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6396 = _T_5 ? offset_215 : _GEN_5359; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6397 = _T_5 ? offset_216 : _GEN_5360; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6398 = _T_5 ? offset_217 : _GEN_5361; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6399 = _T_5 ? offset_218 : _GEN_5362; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6400 = _T_5 ? offset_219 : _GEN_5363; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6401 = _T_5 ? offset_220 : _GEN_5364; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6402 = _T_5 ? offset_221 : _GEN_5365; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6403 = _T_5 ? offset_222 : _GEN_5366; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6404 = _T_5 ? offset_223 : _GEN_5367; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6405 = _T_5 ? offset_224 : _GEN_5368; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6406 = _T_5 ? offset_225 : _GEN_5369; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6407 = _T_5 ? offset_226 : _GEN_5370; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6408 = _T_5 ? offset_227 : _GEN_5371; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6409 = _T_5 ? offset_228 : _GEN_5372; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6410 = _T_5 ? offset_229 : _GEN_5373; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6411 = _T_5 ? offset_230 : _GEN_5374; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6412 = _T_5 ? offset_231 : _GEN_5375; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6413 = _T_5 ? offset_232 : _GEN_5376; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6414 = _T_5 ? offset_233 : _GEN_5377; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6415 = _T_5 ? offset_234 : _GEN_5378; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6416 = _T_5 ? offset_235 : _GEN_5379; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6417 = _T_5 ? offset_236 : _GEN_5380; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6418 = _T_5 ? offset_237 : _GEN_5381; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6419 = _T_5 ? offset_238 : _GEN_5382; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6420 = _T_5 ? offset_239 : _GEN_5383; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6421 = _T_5 ? offset_240 : _GEN_5384; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6422 = _T_5 ? offset_241 : _GEN_5385; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6423 = _T_5 ? offset_242 : _GEN_5386; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6424 = _T_5 ? offset_243 : _GEN_5387; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6425 = _T_5 ? offset_244 : _GEN_5388; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6426 = _T_5 ? offset_245 : _GEN_5389; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6427 = _T_5 ? offset_246 : _GEN_5390; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6428 = _T_5 ? offset_247 : _GEN_5391; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6429 = _T_5 ? offset_248 : _GEN_5392; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6430 = _T_5 ? offset_249 : _GEN_5393; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6431 = _T_5 ? offset_250 : _GEN_5394; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6432 = _T_5 ? offset_251 : _GEN_5395; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6433 = _T_5 ? offset_252 : _GEN_5396; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6434 = _T_5 ? offset_253 : _GEN_5397; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6435 = _T_5 ? offset_254 : _GEN_5398; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_6436 = _T_5 ? offset_255 : _GEN_5399; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [2:0] _GEN_6437 = _T_4 ? 3'h4 : _GEN_5401; // @[Conditional.scala 39:67 Dcache.scala 170:15]
  wire [31:0] _GEN_6438 = _T_4 ? 32'h0 : _GEN_5402; // @[Conditional.scala 39:67]
  wire  _GEN_6442 = _T_4 ? 1'h0 : _T_5 & _GEN_3348; // @[Conditional.scala 39:67]
  wire  _GEN_6444 = _T_4 ? cache_fill : _GEN_5408; // @[Conditional.scala 39:67 Dcache.scala 116:28]
  wire  _GEN_6445 = _T_4 ? cache_wen : _GEN_5409; // @[Conditional.scala 39:67 Dcache.scala 117:28]
  wire [127:0] _GEN_6446 = _T_4 ? cache_wdata : _GEN_5410; // @[Conditional.scala 39:67 Dcache.scala 118:28]
  wire [127:0] _GEN_6447 = _T_4 ? cache_strb : _GEN_5411; // @[Conditional.scala 39:67 Dcache.scala 119:28]
  wire  _GEN_6448 = _T_4 ? data_ready : _GEN_5412; // @[Conditional.scala 39:67 Dcache.scala 46:28]
  wire  _GEN_6449 = _T_4 ? valid_0 : _GEN_5413; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6450 = _T_4 ? valid_1 : _GEN_5414; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6451 = _T_4 ? valid_2 : _GEN_5415; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6452 = _T_4 ? valid_3 : _GEN_5416; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6453 = _T_4 ? valid_4 : _GEN_5417; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6454 = _T_4 ? valid_5 : _GEN_5418; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6455 = _T_4 ? valid_6 : _GEN_5419; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6456 = _T_4 ? valid_7 : _GEN_5420; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6457 = _T_4 ? valid_8 : _GEN_5421; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6458 = _T_4 ? valid_9 : _GEN_5422; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6459 = _T_4 ? valid_10 : _GEN_5423; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6460 = _T_4 ? valid_11 : _GEN_5424; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6461 = _T_4 ? valid_12 : _GEN_5425; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6462 = _T_4 ? valid_13 : _GEN_5426; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6463 = _T_4 ? valid_14 : _GEN_5427; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6464 = _T_4 ? valid_15 : _GEN_5428; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6465 = _T_4 ? valid_16 : _GEN_5429; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6466 = _T_4 ? valid_17 : _GEN_5430; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6467 = _T_4 ? valid_18 : _GEN_5431; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6468 = _T_4 ? valid_19 : _GEN_5432; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6469 = _T_4 ? valid_20 : _GEN_5433; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6470 = _T_4 ? valid_21 : _GEN_5434; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6471 = _T_4 ? valid_22 : _GEN_5435; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6472 = _T_4 ? valid_23 : _GEN_5436; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6473 = _T_4 ? valid_24 : _GEN_5437; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6474 = _T_4 ? valid_25 : _GEN_5438; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6475 = _T_4 ? valid_26 : _GEN_5439; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6476 = _T_4 ? valid_27 : _GEN_5440; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6477 = _T_4 ? valid_28 : _GEN_5441; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6478 = _T_4 ? valid_29 : _GEN_5442; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6479 = _T_4 ? valid_30 : _GEN_5443; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6480 = _T_4 ? valid_31 : _GEN_5444; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6481 = _T_4 ? valid_32 : _GEN_5445; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6482 = _T_4 ? valid_33 : _GEN_5446; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6483 = _T_4 ? valid_34 : _GEN_5447; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6484 = _T_4 ? valid_35 : _GEN_5448; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6485 = _T_4 ? valid_36 : _GEN_5449; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6486 = _T_4 ? valid_37 : _GEN_5450; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6487 = _T_4 ? valid_38 : _GEN_5451; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6488 = _T_4 ? valid_39 : _GEN_5452; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6489 = _T_4 ? valid_40 : _GEN_5453; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6490 = _T_4 ? valid_41 : _GEN_5454; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6491 = _T_4 ? valid_42 : _GEN_5455; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6492 = _T_4 ? valid_43 : _GEN_5456; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6493 = _T_4 ? valid_44 : _GEN_5457; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6494 = _T_4 ? valid_45 : _GEN_5458; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6495 = _T_4 ? valid_46 : _GEN_5459; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6496 = _T_4 ? valid_47 : _GEN_5460; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6497 = _T_4 ? valid_48 : _GEN_5461; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6498 = _T_4 ? valid_49 : _GEN_5462; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6499 = _T_4 ? valid_50 : _GEN_5463; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6500 = _T_4 ? valid_51 : _GEN_5464; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6501 = _T_4 ? valid_52 : _GEN_5465; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6502 = _T_4 ? valid_53 : _GEN_5466; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6503 = _T_4 ? valid_54 : _GEN_5467; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6504 = _T_4 ? valid_55 : _GEN_5468; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6505 = _T_4 ? valid_56 : _GEN_5469; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6506 = _T_4 ? valid_57 : _GEN_5470; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6507 = _T_4 ? valid_58 : _GEN_5471; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6508 = _T_4 ? valid_59 : _GEN_5472; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6509 = _T_4 ? valid_60 : _GEN_5473; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6510 = _T_4 ? valid_61 : _GEN_5474; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6511 = _T_4 ? valid_62 : _GEN_5475; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6512 = _T_4 ? valid_63 : _GEN_5476; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6513 = _T_4 ? valid_64 : _GEN_5477; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6514 = _T_4 ? valid_65 : _GEN_5478; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6515 = _T_4 ? valid_66 : _GEN_5479; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6516 = _T_4 ? valid_67 : _GEN_5480; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6517 = _T_4 ? valid_68 : _GEN_5481; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6518 = _T_4 ? valid_69 : _GEN_5482; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6519 = _T_4 ? valid_70 : _GEN_5483; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6520 = _T_4 ? valid_71 : _GEN_5484; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6521 = _T_4 ? valid_72 : _GEN_5485; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6522 = _T_4 ? valid_73 : _GEN_5486; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6523 = _T_4 ? valid_74 : _GEN_5487; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6524 = _T_4 ? valid_75 : _GEN_5488; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6525 = _T_4 ? valid_76 : _GEN_5489; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6526 = _T_4 ? valid_77 : _GEN_5490; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6527 = _T_4 ? valid_78 : _GEN_5491; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6528 = _T_4 ? valid_79 : _GEN_5492; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6529 = _T_4 ? valid_80 : _GEN_5493; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6530 = _T_4 ? valid_81 : _GEN_5494; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6531 = _T_4 ? valid_82 : _GEN_5495; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6532 = _T_4 ? valid_83 : _GEN_5496; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6533 = _T_4 ? valid_84 : _GEN_5497; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6534 = _T_4 ? valid_85 : _GEN_5498; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6535 = _T_4 ? valid_86 : _GEN_5499; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6536 = _T_4 ? valid_87 : _GEN_5500; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6537 = _T_4 ? valid_88 : _GEN_5501; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6538 = _T_4 ? valid_89 : _GEN_5502; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6539 = _T_4 ? valid_90 : _GEN_5503; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6540 = _T_4 ? valid_91 : _GEN_5504; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6541 = _T_4 ? valid_92 : _GEN_5505; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6542 = _T_4 ? valid_93 : _GEN_5506; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6543 = _T_4 ? valid_94 : _GEN_5507; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6544 = _T_4 ? valid_95 : _GEN_5508; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6545 = _T_4 ? valid_96 : _GEN_5509; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6546 = _T_4 ? valid_97 : _GEN_5510; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6547 = _T_4 ? valid_98 : _GEN_5511; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6548 = _T_4 ? valid_99 : _GEN_5512; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6549 = _T_4 ? valid_100 : _GEN_5513; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6550 = _T_4 ? valid_101 : _GEN_5514; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6551 = _T_4 ? valid_102 : _GEN_5515; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6552 = _T_4 ? valid_103 : _GEN_5516; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6553 = _T_4 ? valid_104 : _GEN_5517; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6554 = _T_4 ? valid_105 : _GEN_5518; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6555 = _T_4 ? valid_106 : _GEN_5519; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6556 = _T_4 ? valid_107 : _GEN_5520; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6557 = _T_4 ? valid_108 : _GEN_5521; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6558 = _T_4 ? valid_109 : _GEN_5522; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6559 = _T_4 ? valid_110 : _GEN_5523; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6560 = _T_4 ? valid_111 : _GEN_5524; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6561 = _T_4 ? valid_112 : _GEN_5525; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6562 = _T_4 ? valid_113 : _GEN_5526; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6563 = _T_4 ? valid_114 : _GEN_5527; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6564 = _T_4 ? valid_115 : _GEN_5528; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6565 = _T_4 ? valid_116 : _GEN_5529; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6566 = _T_4 ? valid_117 : _GEN_5530; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6567 = _T_4 ? valid_118 : _GEN_5531; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6568 = _T_4 ? valid_119 : _GEN_5532; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6569 = _T_4 ? valid_120 : _GEN_5533; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6570 = _T_4 ? valid_121 : _GEN_5534; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6571 = _T_4 ? valid_122 : _GEN_5535; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6572 = _T_4 ? valid_123 : _GEN_5536; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6573 = _T_4 ? valid_124 : _GEN_5537; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6574 = _T_4 ? valid_125 : _GEN_5538; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6575 = _T_4 ? valid_126 : _GEN_5539; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6576 = _T_4 ? valid_127 : _GEN_5540; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6577 = _T_4 ? valid_128 : _GEN_5541; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6578 = _T_4 ? valid_129 : _GEN_5542; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6579 = _T_4 ? valid_130 : _GEN_5543; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6580 = _T_4 ? valid_131 : _GEN_5544; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6581 = _T_4 ? valid_132 : _GEN_5545; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6582 = _T_4 ? valid_133 : _GEN_5546; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6583 = _T_4 ? valid_134 : _GEN_5547; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6584 = _T_4 ? valid_135 : _GEN_5548; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6585 = _T_4 ? valid_136 : _GEN_5549; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6586 = _T_4 ? valid_137 : _GEN_5550; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6587 = _T_4 ? valid_138 : _GEN_5551; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6588 = _T_4 ? valid_139 : _GEN_5552; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6589 = _T_4 ? valid_140 : _GEN_5553; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6590 = _T_4 ? valid_141 : _GEN_5554; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6591 = _T_4 ? valid_142 : _GEN_5555; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6592 = _T_4 ? valid_143 : _GEN_5556; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6593 = _T_4 ? valid_144 : _GEN_5557; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6594 = _T_4 ? valid_145 : _GEN_5558; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6595 = _T_4 ? valid_146 : _GEN_5559; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6596 = _T_4 ? valid_147 : _GEN_5560; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6597 = _T_4 ? valid_148 : _GEN_5561; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6598 = _T_4 ? valid_149 : _GEN_5562; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6599 = _T_4 ? valid_150 : _GEN_5563; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6600 = _T_4 ? valid_151 : _GEN_5564; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6601 = _T_4 ? valid_152 : _GEN_5565; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6602 = _T_4 ? valid_153 : _GEN_5566; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6603 = _T_4 ? valid_154 : _GEN_5567; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6604 = _T_4 ? valid_155 : _GEN_5568; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6605 = _T_4 ? valid_156 : _GEN_5569; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6606 = _T_4 ? valid_157 : _GEN_5570; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6607 = _T_4 ? valid_158 : _GEN_5571; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6608 = _T_4 ? valid_159 : _GEN_5572; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6609 = _T_4 ? valid_160 : _GEN_5573; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6610 = _T_4 ? valid_161 : _GEN_5574; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6611 = _T_4 ? valid_162 : _GEN_5575; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6612 = _T_4 ? valid_163 : _GEN_5576; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6613 = _T_4 ? valid_164 : _GEN_5577; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6614 = _T_4 ? valid_165 : _GEN_5578; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6615 = _T_4 ? valid_166 : _GEN_5579; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6616 = _T_4 ? valid_167 : _GEN_5580; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6617 = _T_4 ? valid_168 : _GEN_5581; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6618 = _T_4 ? valid_169 : _GEN_5582; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6619 = _T_4 ? valid_170 : _GEN_5583; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6620 = _T_4 ? valid_171 : _GEN_5584; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6621 = _T_4 ? valid_172 : _GEN_5585; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6622 = _T_4 ? valid_173 : _GEN_5586; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6623 = _T_4 ? valid_174 : _GEN_5587; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6624 = _T_4 ? valid_175 : _GEN_5588; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6625 = _T_4 ? valid_176 : _GEN_5589; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6626 = _T_4 ? valid_177 : _GEN_5590; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6627 = _T_4 ? valid_178 : _GEN_5591; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6628 = _T_4 ? valid_179 : _GEN_5592; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6629 = _T_4 ? valid_180 : _GEN_5593; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6630 = _T_4 ? valid_181 : _GEN_5594; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6631 = _T_4 ? valid_182 : _GEN_5595; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6632 = _T_4 ? valid_183 : _GEN_5596; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6633 = _T_4 ? valid_184 : _GEN_5597; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6634 = _T_4 ? valid_185 : _GEN_5598; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6635 = _T_4 ? valid_186 : _GEN_5599; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6636 = _T_4 ? valid_187 : _GEN_5600; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6637 = _T_4 ? valid_188 : _GEN_5601; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6638 = _T_4 ? valid_189 : _GEN_5602; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6639 = _T_4 ? valid_190 : _GEN_5603; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6640 = _T_4 ? valid_191 : _GEN_5604; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6641 = _T_4 ? valid_192 : _GEN_5605; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6642 = _T_4 ? valid_193 : _GEN_5606; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6643 = _T_4 ? valid_194 : _GEN_5607; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6644 = _T_4 ? valid_195 : _GEN_5608; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6645 = _T_4 ? valid_196 : _GEN_5609; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6646 = _T_4 ? valid_197 : _GEN_5610; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6647 = _T_4 ? valid_198 : _GEN_5611; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6648 = _T_4 ? valid_199 : _GEN_5612; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6649 = _T_4 ? valid_200 : _GEN_5613; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6650 = _T_4 ? valid_201 : _GEN_5614; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6651 = _T_4 ? valid_202 : _GEN_5615; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6652 = _T_4 ? valid_203 : _GEN_5616; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6653 = _T_4 ? valid_204 : _GEN_5617; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6654 = _T_4 ? valid_205 : _GEN_5618; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6655 = _T_4 ? valid_206 : _GEN_5619; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6656 = _T_4 ? valid_207 : _GEN_5620; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6657 = _T_4 ? valid_208 : _GEN_5621; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6658 = _T_4 ? valid_209 : _GEN_5622; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6659 = _T_4 ? valid_210 : _GEN_5623; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6660 = _T_4 ? valid_211 : _GEN_5624; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6661 = _T_4 ? valid_212 : _GEN_5625; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6662 = _T_4 ? valid_213 : _GEN_5626; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6663 = _T_4 ? valid_214 : _GEN_5627; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6664 = _T_4 ? valid_215 : _GEN_5628; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6665 = _T_4 ? valid_216 : _GEN_5629; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6666 = _T_4 ? valid_217 : _GEN_5630; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6667 = _T_4 ? valid_218 : _GEN_5631; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6668 = _T_4 ? valid_219 : _GEN_5632; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6669 = _T_4 ? valid_220 : _GEN_5633; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6670 = _T_4 ? valid_221 : _GEN_5634; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6671 = _T_4 ? valid_222 : _GEN_5635; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6672 = _T_4 ? valid_223 : _GEN_5636; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6673 = _T_4 ? valid_224 : _GEN_5637; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6674 = _T_4 ? valid_225 : _GEN_5638; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6675 = _T_4 ? valid_226 : _GEN_5639; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6676 = _T_4 ? valid_227 : _GEN_5640; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6677 = _T_4 ? valid_228 : _GEN_5641; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6678 = _T_4 ? valid_229 : _GEN_5642; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6679 = _T_4 ? valid_230 : _GEN_5643; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6680 = _T_4 ? valid_231 : _GEN_5644; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6681 = _T_4 ? valid_232 : _GEN_5645; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6682 = _T_4 ? valid_233 : _GEN_5646; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6683 = _T_4 ? valid_234 : _GEN_5647; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6684 = _T_4 ? valid_235 : _GEN_5648; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6685 = _T_4 ? valid_236 : _GEN_5649; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6686 = _T_4 ? valid_237 : _GEN_5650; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6687 = _T_4 ? valid_238 : _GEN_5651; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6688 = _T_4 ? valid_239 : _GEN_5652; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6689 = _T_4 ? valid_240 : _GEN_5653; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6690 = _T_4 ? valid_241 : _GEN_5654; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6691 = _T_4 ? valid_242 : _GEN_5655; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6692 = _T_4 ? valid_243 : _GEN_5656; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6693 = _T_4 ? valid_244 : _GEN_5657; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6694 = _T_4 ? valid_245 : _GEN_5658; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6695 = _T_4 ? valid_246 : _GEN_5659; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6696 = _T_4 ? valid_247 : _GEN_5660; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6697 = _T_4 ? valid_248 : _GEN_5661; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6698 = _T_4 ? valid_249 : _GEN_5662; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6699 = _T_4 ? valid_250 : _GEN_5663; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6700 = _T_4 ? valid_251 : _GEN_5664; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6701 = _T_4 ? valid_252 : _GEN_5665; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6702 = _T_4 ? valid_253 : _GEN_5666; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6703 = _T_4 ? valid_254 : _GEN_5667; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire  _GEN_6704 = _T_4 ? valid_255 : _GEN_5668; // @[Conditional.scala 39:67 Dcache.scala 17:24]
  wire [19:0] _GEN_6705 = _T_4 ? tag_0 : _GEN_5669; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6706 = _T_4 ? tag_1 : _GEN_5670; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6707 = _T_4 ? tag_2 : _GEN_5671; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6708 = _T_4 ? tag_3 : _GEN_5672; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6709 = _T_4 ? tag_4 : _GEN_5673; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6710 = _T_4 ? tag_5 : _GEN_5674; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6711 = _T_4 ? tag_6 : _GEN_5675; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6712 = _T_4 ? tag_7 : _GEN_5676; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6713 = _T_4 ? tag_8 : _GEN_5677; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6714 = _T_4 ? tag_9 : _GEN_5678; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6715 = _T_4 ? tag_10 : _GEN_5679; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6716 = _T_4 ? tag_11 : _GEN_5680; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6717 = _T_4 ? tag_12 : _GEN_5681; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6718 = _T_4 ? tag_13 : _GEN_5682; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6719 = _T_4 ? tag_14 : _GEN_5683; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6720 = _T_4 ? tag_15 : _GEN_5684; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6721 = _T_4 ? tag_16 : _GEN_5685; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6722 = _T_4 ? tag_17 : _GEN_5686; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6723 = _T_4 ? tag_18 : _GEN_5687; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6724 = _T_4 ? tag_19 : _GEN_5688; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6725 = _T_4 ? tag_20 : _GEN_5689; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6726 = _T_4 ? tag_21 : _GEN_5690; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6727 = _T_4 ? tag_22 : _GEN_5691; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6728 = _T_4 ? tag_23 : _GEN_5692; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6729 = _T_4 ? tag_24 : _GEN_5693; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6730 = _T_4 ? tag_25 : _GEN_5694; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6731 = _T_4 ? tag_26 : _GEN_5695; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6732 = _T_4 ? tag_27 : _GEN_5696; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6733 = _T_4 ? tag_28 : _GEN_5697; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6734 = _T_4 ? tag_29 : _GEN_5698; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6735 = _T_4 ? tag_30 : _GEN_5699; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6736 = _T_4 ? tag_31 : _GEN_5700; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6737 = _T_4 ? tag_32 : _GEN_5701; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6738 = _T_4 ? tag_33 : _GEN_5702; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6739 = _T_4 ? tag_34 : _GEN_5703; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6740 = _T_4 ? tag_35 : _GEN_5704; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6741 = _T_4 ? tag_36 : _GEN_5705; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6742 = _T_4 ? tag_37 : _GEN_5706; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6743 = _T_4 ? tag_38 : _GEN_5707; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6744 = _T_4 ? tag_39 : _GEN_5708; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6745 = _T_4 ? tag_40 : _GEN_5709; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6746 = _T_4 ? tag_41 : _GEN_5710; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6747 = _T_4 ? tag_42 : _GEN_5711; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6748 = _T_4 ? tag_43 : _GEN_5712; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6749 = _T_4 ? tag_44 : _GEN_5713; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6750 = _T_4 ? tag_45 : _GEN_5714; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6751 = _T_4 ? tag_46 : _GEN_5715; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6752 = _T_4 ? tag_47 : _GEN_5716; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6753 = _T_4 ? tag_48 : _GEN_5717; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6754 = _T_4 ? tag_49 : _GEN_5718; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6755 = _T_4 ? tag_50 : _GEN_5719; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6756 = _T_4 ? tag_51 : _GEN_5720; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6757 = _T_4 ? tag_52 : _GEN_5721; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6758 = _T_4 ? tag_53 : _GEN_5722; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6759 = _T_4 ? tag_54 : _GEN_5723; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6760 = _T_4 ? tag_55 : _GEN_5724; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6761 = _T_4 ? tag_56 : _GEN_5725; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6762 = _T_4 ? tag_57 : _GEN_5726; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6763 = _T_4 ? tag_58 : _GEN_5727; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6764 = _T_4 ? tag_59 : _GEN_5728; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6765 = _T_4 ? tag_60 : _GEN_5729; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6766 = _T_4 ? tag_61 : _GEN_5730; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6767 = _T_4 ? tag_62 : _GEN_5731; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6768 = _T_4 ? tag_63 : _GEN_5732; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6769 = _T_4 ? tag_64 : _GEN_5733; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6770 = _T_4 ? tag_65 : _GEN_5734; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6771 = _T_4 ? tag_66 : _GEN_5735; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6772 = _T_4 ? tag_67 : _GEN_5736; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6773 = _T_4 ? tag_68 : _GEN_5737; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6774 = _T_4 ? tag_69 : _GEN_5738; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6775 = _T_4 ? tag_70 : _GEN_5739; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6776 = _T_4 ? tag_71 : _GEN_5740; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6777 = _T_4 ? tag_72 : _GEN_5741; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6778 = _T_4 ? tag_73 : _GEN_5742; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6779 = _T_4 ? tag_74 : _GEN_5743; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6780 = _T_4 ? tag_75 : _GEN_5744; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6781 = _T_4 ? tag_76 : _GEN_5745; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6782 = _T_4 ? tag_77 : _GEN_5746; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6783 = _T_4 ? tag_78 : _GEN_5747; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6784 = _T_4 ? tag_79 : _GEN_5748; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6785 = _T_4 ? tag_80 : _GEN_5749; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6786 = _T_4 ? tag_81 : _GEN_5750; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6787 = _T_4 ? tag_82 : _GEN_5751; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6788 = _T_4 ? tag_83 : _GEN_5752; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6789 = _T_4 ? tag_84 : _GEN_5753; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6790 = _T_4 ? tag_85 : _GEN_5754; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6791 = _T_4 ? tag_86 : _GEN_5755; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6792 = _T_4 ? tag_87 : _GEN_5756; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6793 = _T_4 ? tag_88 : _GEN_5757; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6794 = _T_4 ? tag_89 : _GEN_5758; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6795 = _T_4 ? tag_90 : _GEN_5759; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6796 = _T_4 ? tag_91 : _GEN_5760; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6797 = _T_4 ? tag_92 : _GEN_5761; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6798 = _T_4 ? tag_93 : _GEN_5762; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6799 = _T_4 ? tag_94 : _GEN_5763; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6800 = _T_4 ? tag_95 : _GEN_5764; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6801 = _T_4 ? tag_96 : _GEN_5765; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6802 = _T_4 ? tag_97 : _GEN_5766; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6803 = _T_4 ? tag_98 : _GEN_5767; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6804 = _T_4 ? tag_99 : _GEN_5768; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6805 = _T_4 ? tag_100 : _GEN_5769; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6806 = _T_4 ? tag_101 : _GEN_5770; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6807 = _T_4 ? tag_102 : _GEN_5771; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6808 = _T_4 ? tag_103 : _GEN_5772; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6809 = _T_4 ? tag_104 : _GEN_5773; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6810 = _T_4 ? tag_105 : _GEN_5774; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6811 = _T_4 ? tag_106 : _GEN_5775; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6812 = _T_4 ? tag_107 : _GEN_5776; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6813 = _T_4 ? tag_108 : _GEN_5777; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6814 = _T_4 ? tag_109 : _GEN_5778; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6815 = _T_4 ? tag_110 : _GEN_5779; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6816 = _T_4 ? tag_111 : _GEN_5780; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6817 = _T_4 ? tag_112 : _GEN_5781; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6818 = _T_4 ? tag_113 : _GEN_5782; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6819 = _T_4 ? tag_114 : _GEN_5783; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6820 = _T_4 ? tag_115 : _GEN_5784; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6821 = _T_4 ? tag_116 : _GEN_5785; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6822 = _T_4 ? tag_117 : _GEN_5786; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6823 = _T_4 ? tag_118 : _GEN_5787; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6824 = _T_4 ? tag_119 : _GEN_5788; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6825 = _T_4 ? tag_120 : _GEN_5789; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6826 = _T_4 ? tag_121 : _GEN_5790; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6827 = _T_4 ? tag_122 : _GEN_5791; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6828 = _T_4 ? tag_123 : _GEN_5792; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6829 = _T_4 ? tag_124 : _GEN_5793; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6830 = _T_4 ? tag_125 : _GEN_5794; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6831 = _T_4 ? tag_126 : _GEN_5795; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6832 = _T_4 ? tag_127 : _GEN_5796; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6833 = _T_4 ? tag_128 : _GEN_5797; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6834 = _T_4 ? tag_129 : _GEN_5798; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6835 = _T_4 ? tag_130 : _GEN_5799; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6836 = _T_4 ? tag_131 : _GEN_5800; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6837 = _T_4 ? tag_132 : _GEN_5801; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6838 = _T_4 ? tag_133 : _GEN_5802; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6839 = _T_4 ? tag_134 : _GEN_5803; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6840 = _T_4 ? tag_135 : _GEN_5804; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6841 = _T_4 ? tag_136 : _GEN_5805; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6842 = _T_4 ? tag_137 : _GEN_5806; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6843 = _T_4 ? tag_138 : _GEN_5807; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6844 = _T_4 ? tag_139 : _GEN_5808; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6845 = _T_4 ? tag_140 : _GEN_5809; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6846 = _T_4 ? tag_141 : _GEN_5810; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6847 = _T_4 ? tag_142 : _GEN_5811; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6848 = _T_4 ? tag_143 : _GEN_5812; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6849 = _T_4 ? tag_144 : _GEN_5813; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6850 = _T_4 ? tag_145 : _GEN_5814; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6851 = _T_4 ? tag_146 : _GEN_5815; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6852 = _T_4 ? tag_147 : _GEN_5816; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6853 = _T_4 ? tag_148 : _GEN_5817; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6854 = _T_4 ? tag_149 : _GEN_5818; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6855 = _T_4 ? tag_150 : _GEN_5819; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6856 = _T_4 ? tag_151 : _GEN_5820; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6857 = _T_4 ? tag_152 : _GEN_5821; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6858 = _T_4 ? tag_153 : _GEN_5822; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6859 = _T_4 ? tag_154 : _GEN_5823; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6860 = _T_4 ? tag_155 : _GEN_5824; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6861 = _T_4 ? tag_156 : _GEN_5825; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6862 = _T_4 ? tag_157 : _GEN_5826; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6863 = _T_4 ? tag_158 : _GEN_5827; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6864 = _T_4 ? tag_159 : _GEN_5828; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6865 = _T_4 ? tag_160 : _GEN_5829; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6866 = _T_4 ? tag_161 : _GEN_5830; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6867 = _T_4 ? tag_162 : _GEN_5831; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6868 = _T_4 ? tag_163 : _GEN_5832; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6869 = _T_4 ? tag_164 : _GEN_5833; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6870 = _T_4 ? tag_165 : _GEN_5834; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6871 = _T_4 ? tag_166 : _GEN_5835; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6872 = _T_4 ? tag_167 : _GEN_5836; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6873 = _T_4 ? tag_168 : _GEN_5837; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6874 = _T_4 ? tag_169 : _GEN_5838; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6875 = _T_4 ? tag_170 : _GEN_5839; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6876 = _T_4 ? tag_171 : _GEN_5840; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6877 = _T_4 ? tag_172 : _GEN_5841; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6878 = _T_4 ? tag_173 : _GEN_5842; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6879 = _T_4 ? tag_174 : _GEN_5843; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6880 = _T_4 ? tag_175 : _GEN_5844; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6881 = _T_4 ? tag_176 : _GEN_5845; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6882 = _T_4 ? tag_177 : _GEN_5846; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6883 = _T_4 ? tag_178 : _GEN_5847; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6884 = _T_4 ? tag_179 : _GEN_5848; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6885 = _T_4 ? tag_180 : _GEN_5849; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6886 = _T_4 ? tag_181 : _GEN_5850; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6887 = _T_4 ? tag_182 : _GEN_5851; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6888 = _T_4 ? tag_183 : _GEN_5852; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6889 = _T_4 ? tag_184 : _GEN_5853; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6890 = _T_4 ? tag_185 : _GEN_5854; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6891 = _T_4 ? tag_186 : _GEN_5855; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6892 = _T_4 ? tag_187 : _GEN_5856; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6893 = _T_4 ? tag_188 : _GEN_5857; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6894 = _T_4 ? tag_189 : _GEN_5858; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6895 = _T_4 ? tag_190 : _GEN_5859; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6896 = _T_4 ? tag_191 : _GEN_5860; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6897 = _T_4 ? tag_192 : _GEN_5861; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6898 = _T_4 ? tag_193 : _GEN_5862; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6899 = _T_4 ? tag_194 : _GEN_5863; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6900 = _T_4 ? tag_195 : _GEN_5864; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6901 = _T_4 ? tag_196 : _GEN_5865; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6902 = _T_4 ? tag_197 : _GEN_5866; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6903 = _T_4 ? tag_198 : _GEN_5867; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6904 = _T_4 ? tag_199 : _GEN_5868; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6905 = _T_4 ? tag_200 : _GEN_5869; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6906 = _T_4 ? tag_201 : _GEN_5870; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6907 = _T_4 ? tag_202 : _GEN_5871; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6908 = _T_4 ? tag_203 : _GEN_5872; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6909 = _T_4 ? tag_204 : _GEN_5873; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6910 = _T_4 ? tag_205 : _GEN_5874; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6911 = _T_4 ? tag_206 : _GEN_5875; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6912 = _T_4 ? tag_207 : _GEN_5876; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6913 = _T_4 ? tag_208 : _GEN_5877; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6914 = _T_4 ? tag_209 : _GEN_5878; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6915 = _T_4 ? tag_210 : _GEN_5879; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6916 = _T_4 ? tag_211 : _GEN_5880; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6917 = _T_4 ? tag_212 : _GEN_5881; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6918 = _T_4 ? tag_213 : _GEN_5882; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6919 = _T_4 ? tag_214 : _GEN_5883; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6920 = _T_4 ? tag_215 : _GEN_5884; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6921 = _T_4 ? tag_216 : _GEN_5885; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6922 = _T_4 ? tag_217 : _GEN_5886; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6923 = _T_4 ? tag_218 : _GEN_5887; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6924 = _T_4 ? tag_219 : _GEN_5888; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6925 = _T_4 ? tag_220 : _GEN_5889; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6926 = _T_4 ? tag_221 : _GEN_5890; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6927 = _T_4 ? tag_222 : _GEN_5891; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6928 = _T_4 ? tag_223 : _GEN_5892; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6929 = _T_4 ? tag_224 : _GEN_5893; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6930 = _T_4 ? tag_225 : _GEN_5894; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6931 = _T_4 ? tag_226 : _GEN_5895; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6932 = _T_4 ? tag_227 : _GEN_5896; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6933 = _T_4 ? tag_228 : _GEN_5897; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6934 = _T_4 ? tag_229 : _GEN_5898; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6935 = _T_4 ? tag_230 : _GEN_5899; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6936 = _T_4 ? tag_231 : _GEN_5900; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6937 = _T_4 ? tag_232 : _GEN_5901; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6938 = _T_4 ? tag_233 : _GEN_5902; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6939 = _T_4 ? tag_234 : _GEN_5903; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6940 = _T_4 ? tag_235 : _GEN_5904; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6941 = _T_4 ? tag_236 : _GEN_5905; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6942 = _T_4 ? tag_237 : _GEN_5906; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6943 = _T_4 ? tag_238 : _GEN_5907; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6944 = _T_4 ? tag_239 : _GEN_5908; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6945 = _T_4 ? tag_240 : _GEN_5909; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6946 = _T_4 ? tag_241 : _GEN_5910; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6947 = _T_4 ? tag_242 : _GEN_5911; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6948 = _T_4 ? tag_243 : _GEN_5912; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6949 = _T_4 ? tag_244 : _GEN_5913; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6950 = _T_4 ? tag_245 : _GEN_5914; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6951 = _T_4 ? tag_246 : _GEN_5915; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6952 = _T_4 ? tag_247 : _GEN_5916; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6953 = _T_4 ? tag_248 : _GEN_5917; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6954 = _T_4 ? tag_249 : _GEN_5918; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6955 = _T_4 ? tag_250 : _GEN_5919; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6956 = _T_4 ? tag_251 : _GEN_5920; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6957 = _T_4 ? tag_252 : _GEN_5921; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6958 = _T_4 ? tag_253 : _GEN_5922; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6959 = _T_4 ? tag_254 : _GEN_5923; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire [19:0] _GEN_6960 = _T_4 ? tag_255 : _GEN_5924; // @[Conditional.scala 39:67 Dcache.scala 16:24]
  wire  _GEN_6961 = _T_4 ? dirty_0 : _GEN_5925; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6962 = _T_4 ? dirty_1 : _GEN_5926; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6963 = _T_4 ? dirty_2 : _GEN_5927; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6964 = _T_4 ? dirty_3 : _GEN_5928; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6965 = _T_4 ? dirty_4 : _GEN_5929; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6966 = _T_4 ? dirty_5 : _GEN_5930; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6967 = _T_4 ? dirty_6 : _GEN_5931; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6968 = _T_4 ? dirty_7 : _GEN_5932; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6969 = _T_4 ? dirty_8 : _GEN_5933; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6970 = _T_4 ? dirty_9 : _GEN_5934; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6971 = _T_4 ? dirty_10 : _GEN_5935; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6972 = _T_4 ? dirty_11 : _GEN_5936; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6973 = _T_4 ? dirty_12 : _GEN_5937; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6974 = _T_4 ? dirty_13 : _GEN_5938; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6975 = _T_4 ? dirty_14 : _GEN_5939; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6976 = _T_4 ? dirty_15 : _GEN_5940; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6977 = _T_4 ? dirty_16 : _GEN_5941; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6978 = _T_4 ? dirty_17 : _GEN_5942; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6979 = _T_4 ? dirty_18 : _GEN_5943; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6980 = _T_4 ? dirty_19 : _GEN_5944; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6981 = _T_4 ? dirty_20 : _GEN_5945; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6982 = _T_4 ? dirty_21 : _GEN_5946; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6983 = _T_4 ? dirty_22 : _GEN_5947; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6984 = _T_4 ? dirty_23 : _GEN_5948; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6985 = _T_4 ? dirty_24 : _GEN_5949; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6986 = _T_4 ? dirty_25 : _GEN_5950; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6987 = _T_4 ? dirty_26 : _GEN_5951; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6988 = _T_4 ? dirty_27 : _GEN_5952; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6989 = _T_4 ? dirty_28 : _GEN_5953; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6990 = _T_4 ? dirty_29 : _GEN_5954; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6991 = _T_4 ? dirty_30 : _GEN_5955; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6992 = _T_4 ? dirty_31 : _GEN_5956; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6993 = _T_4 ? dirty_32 : _GEN_5957; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6994 = _T_4 ? dirty_33 : _GEN_5958; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6995 = _T_4 ? dirty_34 : _GEN_5959; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6996 = _T_4 ? dirty_35 : _GEN_5960; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6997 = _T_4 ? dirty_36 : _GEN_5961; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6998 = _T_4 ? dirty_37 : _GEN_5962; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_6999 = _T_4 ? dirty_38 : _GEN_5963; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7000 = _T_4 ? dirty_39 : _GEN_5964; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7001 = _T_4 ? dirty_40 : _GEN_5965; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7002 = _T_4 ? dirty_41 : _GEN_5966; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7003 = _T_4 ? dirty_42 : _GEN_5967; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7004 = _T_4 ? dirty_43 : _GEN_5968; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7005 = _T_4 ? dirty_44 : _GEN_5969; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7006 = _T_4 ? dirty_45 : _GEN_5970; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7007 = _T_4 ? dirty_46 : _GEN_5971; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7008 = _T_4 ? dirty_47 : _GEN_5972; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7009 = _T_4 ? dirty_48 : _GEN_5973; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7010 = _T_4 ? dirty_49 : _GEN_5974; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7011 = _T_4 ? dirty_50 : _GEN_5975; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7012 = _T_4 ? dirty_51 : _GEN_5976; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7013 = _T_4 ? dirty_52 : _GEN_5977; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7014 = _T_4 ? dirty_53 : _GEN_5978; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7015 = _T_4 ? dirty_54 : _GEN_5979; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7016 = _T_4 ? dirty_55 : _GEN_5980; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7017 = _T_4 ? dirty_56 : _GEN_5981; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7018 = _T_4 ? dirty_57 : _GEN_5982; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7019 = _T_4 ? dirty_58 : _GEN_5983; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7020 = _T_4 ? dirty_59 : _GEN_5984; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7021 = _T_4 ? dirty_60 : _GEN_5985; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7022 = _T_4 ? dirty_61 : _GEN_5986; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7023 = _T_4 ? dirty_62 : _GEN_5987; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7024 = _T_4 ? dirty_63 : _GEN_5988; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7025 = _T_4 ? dirty_64 : _GEN_5989; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7026 = _T_4 ? dirty_65 : _GEN_5990; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7027 = _T_4 ? dirty_66 : _GEN_5991; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7028 = _T_4 ? dirty_67 : _GEN_5992; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7029 = _T_4 ? dirty_68 : _GEN_5993; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7030 = _T_4 ? dirty_69 : _GEN_5994; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7031 = _T_4 ? dirty_70 : _GEN_5995; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7032 = _T_4 ? dirty_71 : _GEN_5996; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7033 = _T_4 ? dirty_72 : _GEN_5997; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7034 = _T_4 ? dirty_73 : _GEN_5998; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7035 = _T_4 ? dirty_74 : _GEN_5999; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7036 = _T_4 ? dirty_75 : _GEN_6000; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7037 = _T_4 ? dirty_76 : _GEN_6001; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7038 = _T_4 ? dirty_77 : _GEN_6002; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7039 = _T_4 ? dirty_78 : _GEN_6003; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7040 = _T_4 ? dirty_79 : _GEN_6004; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7041 = _T_4 ? dirty_80 : _GEN_6005; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7042 = _T_4 ? dirty_81 : _GEN_6006; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7043 = _T_4 ? dirty_82 : _GEN_6007; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7044 = _T_4 ? dirty_83 : _GEN_6008; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7045 = _T_4 ? dirty_84 : _GEN_6009; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7046 = _T_4 ? dirty_85 : _GEN_6010; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7047 = _T_4 ? dirty_86 : _GEN_6011; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7048 = _T_4 ? dirty_87 : _GEN_6012; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7049 = _T_4 ? dirty_88 : _GEN_6013; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7050 = _T_4 ? dirty_89 : _GEN_6014; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7051 = _T_4 ? dirty_90 : _GEN_6015; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7052 = _T_4 ? dirty_91 : _GEN_6016; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7053 = _T_4 ? dirty_92 : _GEN_6017; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7054 = _T_4 ? dirty_93 : _GEN_6018; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7055 = _T_4 ? dirty_94 : _GEN_6019; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7056 = _T_4 ? dirty_95 : _GEN_6020; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7057 = _T_4 ? dirty_96 : _GEN_6021; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7058 = _T_4 ? dirty_97 : _GEN_6022; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7059 = _T_4 ? dirty_98 : _GEN_6023; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7060 = _T_4 ? dirty_99 : _GEN_6024; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7061 = _T_4 ? dirty_100 : _GEN_6025; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7062 = _T_4 ? dirty_101 : _GEN_6026; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7063 = _T_4 ? dirty_102 : _GEN_6027; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7064 = _T_4 ? dirty_103 : _GEN_6028; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7065 = _T_4 ? dirty_104 : _GEN_6029; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7066 = _T_4 ? dirty_105 : _GEN_6030; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7067 = _T_4 ? dirty_106 : _GEN_6031; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7068 = _T_4 ? dirty_107 : _GEN_6032; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7069 = _T_4 ? dirty_108 : _GEN_6033; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7070 = _T_4 ? dirty_109 : _GEN_6034; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7071 = _T_4 ? dirty_110 : _GEN_6035; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7072 = _T_4 ? dirty_111 : _GEN_6036; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7073 = _T_4 ? dirty_112 : _GEN_6037; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7074 = _T_4 ? dirty_113 : _GEN_6038; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7075 = _T_4 ? dirty_114 : _GEN_6039; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7076 = _T_4 ? dirty_115 : _GEN_6040; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7077 = _T_4 ? dirty_116 : _GEN_6041; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7078 = _T_4 ? dirty_117 : _GEN_6042; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7079 = _T_4 ? dirty_118 : _GEN_6043; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7080 = _T_4 ? dirty_119 : _GEN_6044; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7081 = _T_4 ? dirty_120 : _GEN_6045; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7082 = _T_4 ? dirty_121 : _GEN_6046; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7083 = _T_4 ? dirty_122 : _GEN_6047; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7084 = _T_4 ? dirty_123 : _GEN_6048; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7085 = _T_4 ? dirty_124 : _GEN_6049; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7086 = _T_4 ? dirty_125 : _GEN_6050; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7087 = _T_4 ? dirty_126 : _GEN_6051; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7088 = _T_4 ? dirty_127 : _GEN_6052; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7089 = _T_4 ? dirty_128 : _GEN_6053; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7090 = _T_4 ? dirty_129 : _GEN_6054; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7091 = _T_4 ? dirty_130 : _GEN_6055; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7092 = _T_4 ? dirty_131 : _GEN_6056; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7093 = _T_4 ? dirty_132 : _GEN_6057; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7094 = _T_4 ? dirty_133 : _GEN_6058; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7095 = _T_4 ? dirty_134 : _GEN_6059; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7096 = _T_4 ? dirty_135 : _GEN_6060; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7097 = _T_4 ? dirty_136 : _GEN_6061; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7098 = _T_4 ? dirty_137 : _GEN_6062; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7099 = _T_4 ? dirty_138 : _GEN_6063; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7100 = _T_4 ? dirty_139 : _GEN_6064; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7101 = _T_4 ? dirty_140 : _GEN_6065; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7102 = _T_4 ? dirty_141 : _GEN_6066; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7103 = _T_4 ? dirty_142 : _GEN_6067; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7104 = _T_4 ? dirty_143 : _GEN_6068; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7105 = _T_4 ? dirty_144 : _GEN_6069; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7106 = _T_4 ? dirty_145 : _GEN_6070; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7107 = _T_4 ? dirty_146 : _GEN_6071; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7108 = _T_4 ? dirty_147 : _GEN_6072; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7109 = _T_4 ? dirty_148 : _GEN_6073; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7110 = _T_4 ? dirty_149 : _GEN_6074; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7111 = _T_4 ? dirty_150 : _GEN_6075; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7112 = _T_4 ? dirty_151 : _GEN_6076; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7113 = _T_4 ? dirty_152 : _GEN_6077; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7114 = _T_4 ? dirty_153 : _GEN_6078; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7115 = _T_4 ? dirty_154 : _GEN_6079; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7116 = _T_4 ? dirty_155 : _GEN_6080; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7117 = _T_4 ? dirty_156 : _GEN_6081; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7118 = _T_4 ? dirty_157 : _GEN_6082; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7119 = _T_4 ? dirty_158 : _GEN_6083; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7120 = _T_4 ? dirty_159 : _GEN_6084; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7121 = _T_4 ? dirty_160 : _GEN_6085; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7122 = _T_4 ? dirty_161 : _GEN_6086; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7123 = _T_4 ? dirty_162 : _GEN_6087; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7124 = _T_4 ? dirty_163 : _GEN_6088; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7125 = _T_4 ? dirty_164 : _GEN_6089; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7126 = _T_4 ? dirty_165 : _GEN_6090; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7127 = _T_4 ? dirty_166 : _GEN_6091; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7128 = _T_4 ? dirty_167 : _GEN_6092; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7129 = _T_4 ? dirty_168 : _GEN_6093; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7130 = _T_4 ? dirty_169 : _GEN_6094; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7131 = _T_4 ? dirty_170 : _GEN_6095; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7132 = _T_4 ? dirty_171 : _GEN_6096; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7133 = _T_4 ? dirty_172 : _GEN_6097; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7134 = _T_4 ? dirty_173 : _GEN_6098; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7135 = _T_4 ? dirty_174 : _GEN_6099; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7136 = _T_4 ? dirty_175 : _GEN_6100; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7137 = _T_4 ? dirty_176 : _GEN_6101; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7138 = _T_4 ? dirty_177 : _GEN_6102; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7139 = _T_4 ? dirty_178 : _GEN_6103; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7140 = _T_4 ? dirty_179 : _GEN_6104; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7141 = _T_4 ? dirty_180 : _GEN_6105; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7142 = _T_4 ? dirty_181 : _GEN_6106; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7143 = _T_4 ? dirty_182 : _GEN_6107; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7144 = _T_4 ? dirty_183 : _GEN_6108; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7145 = _T_4 ? dirty_184 : _GEN_6109; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7146 = _T_4 ? dirty_185 : _GEN_6110; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7147 = _T_4 ? dirty_186 : _GEN_6111; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7148 = _T_4 ? dirty_187 : _GEN_6112; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7149 = _T_4 ? dirty_188 : _GEN_6113; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7150 = _T_4 ? dirty_189 : _GEN_6114; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7151 = _T_4 ? dirty_190 : _GEN_6115; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7152 = _T_4 ? dirty_191 : _GEN_6116; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7153 = _T_4 ? dirty_192 : _GEN_6117; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7154 = _T_4 ? dirty_193 : _GEN_6118; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7155 = _T_4 ? dirty_194 : _GEN_6119; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7156 = _T_4 ? dirty_195 : _GEN_6120; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7157 = _T_4 ? dirty_196 : _GEN_6121; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7158 = _T_4 ? dirty_197 : _GEN_6122; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7159 = _T_4 ? dirty_198 : _GEN_6123; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7160 = _T_4 ? dirty_199 : _GEN_6124; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7161 = _T_4 ? dirty_200 : _GEN_6125; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7162 = _T_4 ? dirty_201 : _GEN_6126; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7163 = _T_4 ? dirty_202 : _GEN_6127; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7164 = _T_4 ? dirty_203 : _GEN_6128; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7165 = _T_4 ? dirty_204 : _GEN_6129; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7166 = _T_4 ? dirty_205 : _GEN_6130; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7167 = _T_4 ? dirty_206 : _GEN_6131; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7168 = _T_4 ? dirty_207 : _GEN_6132; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7169 = _T_4 ? dirty_208 : _GEN_6133; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7170 = _T_4 ? dirty_209 : _GEN_6134; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7171 = _T_4 ? dirty_210 : _GEN_6135; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7172 = _T_4 ? dirty_211 : _GEN_6136; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7173 = _T_4 ? dirty_212 : _GEN_6137; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7174 = _T_4 ? dirty_213 : _GEN_6138; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7175 = _T_4 ? dirty_214 : _GEN_6139; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7176 = _T_4 ? dirty_215 : _GEN_6140; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7177 = _T_4 ? dirty_216 : _GEN_6141; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7178 = _T_4 ? dirty_217 : _GEN_6142; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7179 = _T_4 ? dirty_218 : _GEN_6143; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7180 = _T_4 ? dirty_219 : _GEN_6144; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7181 = _T_4 ? dirty_220 : _GEN_6145; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7182 = _T_4 ? dirty_221 : _GEN_6146; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7183 = _T_4 ? dirty_222 : _GEN_6147; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7184 = _T_4 ? dirty_223 : _GEN_6148; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7185 = _T_4 ? dirty_224 : _GEN_6149; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7186 = _T_4 ? dirty_225 : _GEN_6150; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7187 = _T_4 ? dirty_226 : _GEN_6151; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7188 = _T_4 ? dirty_227 : _GEN_6152; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7189 = _T_4 ? dirty_228 : _GEN_6153; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7190 = _T_4 ? dirty_229 : _GEN_6154; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7191 = _T_4 ? dirty_230 : _GEN_6155; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7192 = _T_4 ? dirty_231 : _GEN_6156; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7193 = _T_4 ? dirty_232 : _GEN_6157; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7194 = _T_4 ? dirty_233 : _GEN_6158; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7195 = _T_4 ? dirty_234 : _GEN_6159; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7196 = _T_4 ? dirty_235 : _GEN_6160; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7197 = _T_4 ? dirty_236 : _GEN_6161; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7198 = _T_4 ? dirty_237 : _GEN_6162; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7199 = _T_4 ? dirty_238 : _GEN_6163; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7200 = _T_4 ? dirty_239 : _GEN_6164; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7201 = _T_4 ? dirty_240 : _GEN_6165; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7202 = _T_4 ? dirty_241 : _GEN_6166; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7203 = _T_4 ? dirty_242 : _GEN_6167; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7204 = _T_4 ? dirty_243 : _GEN_6168; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7205 = _T_4 ? dirty_244 : _GEN_6169; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7206 = _T_4 ? dirty_245 : _GEN_6170; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7207 = _T_4 ? dirty_246 : _GEN_6171; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7208 = _T_4 ? dirty_247 : _GEN_6172; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7209 = _T_4 ? dirty_248 : _GEN_6173; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7210 = _T_4 ? dirty_249 : _GEN_6174; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7211 = _T_4 ? dirty_250 : _GEN_6175; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7212 = _T_4 ? dirty_251 : _GEN_6176; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7213 = _T_4 ? dirty_252 : _GEN_6177; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7214 = _T_4 ? dirty_253 : _GEN_6178; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7215 = _T_4 ? dirty_254 : _GEN_6179; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire  _GEN_7216 = _T_4 ? dirty_255 : _GEN_6180; // @[Conditional.scala 39:67 Dcache.scala 18:24]
  wire [3:0] _GEN_7217 = _T_4 ? offset_0 : _GEN_6181; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7218 = _T_4 ? offset_1 : _GEN_6182; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7219 = _T_4 ? offset_2 : _GEN_6183; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7220 = _T_4 ? offset_3 : _GEN_6184; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7221 = _T_4 ? offset_4 : _GEN_6185; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7222 = _T_4 ? offset_5 : _GEN_6186; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7223 = _T_4 ? offset_6 : _GEN_6187; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7224 = _T_4 ? offset_7 : _GEN_6188; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7225 = _T_4 ? offset_8 : _GEN_6189; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7226 = _T_4 ? offset_9 : _GEN_6190; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7227 = _T_4 ? offset_10 : _GEN_6191; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7228 = _T_4 ? offset_11 : _GEN_6192; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7229 = _T_4 ? offset_12 : _GEN_6193; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7230 = _T_4 ? offset_13 : _GEN_6194; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7231 = _T_4 ? offset_14 : _GEN_6195; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7232 = _T_4 ? offset_15 : _GEN_6196; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7233 = _T_4 ? offset_16 : _GEN_6197; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7234 = _T_4 ? offset_17 : _GEN_6198; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7235 = _T_4 ? offset_18 : _GEN_6199; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7236 = _T_4 ? offset_19 : _GEN_6200; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7237 = _T_4 ? offset_20 : _GEN_6201; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7238 = _T_4 ? offset_21 : _GEN_6202; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7239 = _T_4 ? offset_22 : _GEN_6203; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7240 = _T_4 ? offset_23 : _GEN_6204; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7241 = _T_4 ? offset_24 : _GEN_6205; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7242 = _T_4 ? offset_25 : _GEN_6206; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7243 = _T_4 ? offset_26 : _GEN_6207; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7244 = _T_4 ? offset_27 : _GEN_6208; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7245 = _T_4 ? offset_28 : _GEN_6209; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7246 = _T_4 ? offset_29 : _GEN_6210; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7247 = _T_4 ? offset_30 : _GEN_6211; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7248 = _T_4 ? offset_31 : _GEN_6212; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7249 = _T_4 ? offset_32 : _GEN_6213; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7250 = _T_4 ? offset_33 : _GEN_6214; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7251 = _T_4 ? offset_34 : _GEN_6215; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7252 = _T_4 ? offset_35 : _GEN_6216; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7253 = _T_4 ? offset_36 : _GEN_6217; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7254 = _T_4 ? offset_37 : _GEN_6218; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7255 = _T_4 ? offset_38 : _GEN_6219; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7256 = _T_4 ? offset_39 : _GEN_6220; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7257 = _T_4 ? offset_40 : _GEN_6221; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7258 = _T_4 ? offset_41 : _GEN_6222; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7259 = _T_4 ? offset_42 : _GEN_6223; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7260 = _T_4 ? offset_43 : _GEN_6224; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7261 = _T_4 ? offset_44 : _GEN_6225; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7262 = _T_4 ? offset_45 : _GEN_6226; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7263 = _T_4 ? offset_46 : _GEN_6227; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7264 = _T_4 ? offset_47 : _GEN_6228; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7265 = _T_4 ? offset_48 : _GEN_6229; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7266 = _T_4 ? offset_49 : _GEN_6230; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7267 = _T_4 ? offset_50 : _GEN_6231; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7268 = _T_4 ? offset_51 : _GEN_6232; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7269 = _T_4 ? offset_52 : _GEN_6233; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7270 = _T_4 ? offset_53 : _GEN_6234; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7271 = _T_4 ? offset_54 : _GEN_6235; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7272 = _T_4 ? offset_55 : _GEN_6236; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7273 = _T_4 ? offset_56 : _GEN_6237; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7274 = _T_4 ? offset_57 : _GEN_6238; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7275 = _T_4 ? offset_58 : _GEN_6239; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7276 = _T_4 ? offset_59 : _GEN_6240; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7277 = _T_4 ? offset_60 : _GEN_6241; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7278 = _T_4 ? offset_61 : _GEN_6242; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7279 = _T_4 ? offset_62 : _GEN_6243; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7280 = _T_4 ? offset_63 : _GEN_6244; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7281 = _T_4 ? offset_64 : _GEN_6245; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7282 = _T_4 ? offset_65 : _GEN_6246; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7283 = _T_4 ? offset_66 : _GEN_6247; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7284 = _T_4 ? offset_67 : _GEN_6248; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7285 = _T_4 ? offset_68 : _GEN_6249; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7286 = _T_4 ? offset_69 : _GEN_6250; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7287 = _T_4 ? offset_70 : _GEN_6251; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7288 = _T_4 ? offset_71 : _GEN_6252; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7289 = _T_4 ? offset_72 : _GEN_6253; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7290 = _T_4 ? offset_73 : _GEN_6254; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7291 = _T_4 ? offset_74 : _GEN_6255; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7292 = _T_4 ? offset_75 : _GEN_6256; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7293 = _T_4 ? offset_76 : _GEN_6257; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7294 = _T_4 ? offset_77 : _GEN_6258; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7295 = _T_4 ? offset_78 : _GEN_6259; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7296 = _T_4 ? offset_79 : _GEN_6260; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7297 = _T_4 ? offset_80 : _GEN_6261; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7298 = _T_4 ? offset_81 : _GEN_6262; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7299 = _T_4 ? offset_82 : _GEN_6263; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7300 = _T_4 ? offset_83 : _GEN_6264; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7301 = _T_4 ? offset_84 : _GEN_6265; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7302 = _T_4 ? offset_85 : _GEN_6266; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7303 = _T_4 ? offset_86 : _GEN_6267; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7304 = _T_4 ? offset_87 : _GEN_6268; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7305 = _T_4 ? offset_88 : _GEN_6269; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7306 = _T_4 ? offset_89 : _GEN_6270; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7307 = _T_4 ? offset_90 : _GEN_6271; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7308 = _T_4 ? offset_91 : _GEN_6272; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7309 = _T_4 ? offset_92 : _GEN_6273; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7310 = _T_4 ? offset_93 : _GEN_6274; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7311 = _T_4 ? offset_94 : _GEN_6275; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7312 = _T_4 ? offset_95 : _GEN_6276; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7313 = _T_4 ? offset_96 : _GEN_6277; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7314 = _T_4 ? offset_97 : _GEN_6278; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7315 = _T_4 ? offset_98 : _GEN_6279; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7316 = _T_4 ? offset_99 : _GEN_6280; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7317 = _T_4 ? offset_100 : _GEN_6281; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7318 = _T_4 ? offset_101 : _GEN_6282; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7319 = _T_4 ? offset_102 : _GEN_6283; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7320 = _T_4 ? offset_103 : _GEN_6284; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7321 = _T_4 ? offset_104 : _GEN_6285; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7322 = _T_4 ? offset_105 : _GEN_6286; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7323 = _T_4 ? offset_106 : _GEN_6287; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7324 = _T_4 ? offset_107 : _GEN_6288; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7325 = _T_4 ? offset_108 : _GEN_6289; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7326 = _T_4 ? offset_109 : _GEN_6290; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7327 = _T_4 ? offset_110 : _GEN_6291; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7328 = _T_4 ? offset_111 : _GEN_6292; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7329 = _T_4 ? offset_112 : _GEN_6293; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7330 = _T_4 ? offset_113 : _GEN_6294; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7331 = _T_4 ? offset_114 : _GEN_6295; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7332 = _T_4 ? offset_115 : _GEN_6296; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7333 = _T_4 ? offset_116 : _GEN_6297; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7334 = _T_4 ? offset_117 : _GEN_6298; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7335 = _T_4 ? offset_118 : _GEN_6299; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7336 = _T_4 ? offset_119 : _GEN_6300; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7337 = _T_4 ? offset_120 : _GEN_6301; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7338 = _T_4 ? offset_121 : _GEN_6302; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7339 = _T_4 ? offset_122 : _GEN_6303; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7340 = _T_4 ? offset_123 : _GEN_6304; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7341 = _T_4 ? offset_124 : _GEN_6305; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7342 = _T_4 ? offset_125 : _GEN_6306; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7343 = _T_4 ? offset_126 : _GEN_6307; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7344 = _T_4 ? offset_127 : _GEN_6308; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7345 = _T_4 ? offset_128 : _GEN_6309; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7346 = _T_4 ? offset_129 : _GEN_6310; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7347 = _T_4 ? offset_130 : _GEN_6311; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7348 = _T_4 ? offset_131 : _GEN_6312; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7349 = _T_4 ? offset_132 : _GEN_6313; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7350 = _T_4 ? offset_133 : _GEN_6314; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7351 = _T_4 ? offset_134 : _GEN_6315; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7352 = _T_4 ? offset_135 : _GEN_6316; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7353 = _T_4 ? offset_136 : _GEN_6317; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7354 = _T_4 ? offset_137 : _GEN_6318; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7355 = _T_4 ? offset_138 : _GEN_6319; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7356 = _T_4 ? offset_139 : _GEN_6320; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7357 = _T_4 ? offset_140 : _GEN_6321; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7358 = _T_4 ? offset_141 : _GEN_6322; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7359 = _T_4 ? offset_142 : _GEN_6323; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7360 = _T_4 ? offset_143 : _GEN_6324; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7361 = _T_4 ? offset_144 : _GEN_6325; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7362 = _T_4 ? offset_145 : _GEN_6326; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7363 = _T_4 ? offset_146 : _GEN_6327; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7364 = _T_4 ? offset_147 : _GEN_6328; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7365 = _T_4 ? offset_148 : _GEN_6329; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7366 = _T_4 ? offset_149 : _GEN_6330; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7367 = _T_4 ? offset_150 : _GEN_6331; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7368 = _T_4 ? offset_151 : _GEN_6332; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7369 = _T_4 ? offset_152 : _GEN_6333; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7370 = _T_4 ? offset_153 : _GEN_6334; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7371 = _T_4 ? offset_154 : _GEN_6335; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7372 = _T_4 ? offset_155 : _GEN_6336; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7373 = _T_4 ? offset_156 : _GEN_6337; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7374 = _T_4 ? offset_157 : _GEN_6338; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7375 = _T_4 ? offset_158 : _GEN_6339; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7376 = _T_4 ? offset_159 : _GEN_6340; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7377 = _T_4 ? offset_160 : _GEN_6341; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7378 = _T_4 ? offset_161 : _GEN_6342; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7379 = _T_4 ? offset_162 : _GEN_6343; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7380 = _T_4 ? offset_163 : _GEN_6344; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7381 = _T_4 ? offset_164 : _GEN_6345; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7382 = _T_4 ? offset_165 : _GEN_6346; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7383 = _T_4 ? offset_166 : _GEN_6347; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7384 = _T_4 ? offset_167 : _GEN_6348; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7385 = _T_4 ? offset_168 : _GEN_6349; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7386 = _T_4 ? offset_169 : _GEN_6350; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7387 = _T_4 ? offset_170 : _GEN_6351; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7388 = _T_4 ? offset_171 : _GEN_6352; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7389 = _T_4 ? offset_172 : _GEN_6353; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7390 = _T_4 ? offset_173 : _GEN_6354; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7391 = _T_4 ? offset_174 : _GEN_6355; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7392 = _T_4 ? offset_175 : _GEN_6356; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7393 = _T_4 ? offset_176 : _GEN_6357; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7394 = _T_4 ? offset_177 : _GEN_6358; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7395 = _T_4 ? offset_178 : _GEN_6359; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7396 = _T_4 ? offset_179 : _GEN_6360; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7397 = _T_4 ? offset_180 : _GEN_6361; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7398 = _T_4 ? offset_181 : _GEN_6362; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7399 = _T_4 ? offset_182 : _GEN_6363; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7400 = _T_4 ? offset_183 : _GEN_6364; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7401 = _T_4 ? offset_184 : _GEN_6365; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7402 = _T_4 ? offset_185 : _GEN_6366; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7403 = _T_4 ? offset_186 : _GEN_6367; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7404 = _T_4 ? offset_187 : _GEN_6368; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7405 = _T_4 ? offset_188 : _GEN_6369; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7406 = _T_4 ? offset_189 : _GEN_6370; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7407 = _T_4 ? offset_190 : _GEN_6371; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7408 = _T_4 ? offset_191 : _GEN_6372; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7409 = _T_4 ? offset_192 : _GEN_6373; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7410 = _T_4 ? offset_193 : _GEN_6374; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7411 = _T_4 ? offset_194 : _GEN_6375; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7412 = _T_4 ? offset_195 : _GEN_6376; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7413 = _T_4 ? offset_196 : _GEN_6377; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7414 = _T_4 ? offset_197 : _GEN_6378; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7415 = _T_4 ? offset_198 : _GEN_6379; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7416 = _T_4 ? offset_199 : _GEN_6380; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7417 = _T_4 ? offset_200 : _GEN_6381; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7418 = _T_4 ? offset_201 : _GEN_6382; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7419 = _T_4 ? offset_202 : _GEN_6383; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7420 = _T_4 ? offset_203 : _GEN_6384; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7421 = _T_4 ? offset_204 : _GEN_6385; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7422 = _T_4 ? offset_205 : _GEN_6386; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7423 = _T_4 ? offset_206 : _GEN_6387; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7424 = _T_4 ? offset_207 : _GEN_6388; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7425 = _T_4 ? offset_208 : _GEN_6389; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7426 = _T_4 ? offset_209 : _GEN_6390; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7427 = _T_4 ? offset_210 : _GEN_6391; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7428 = _T_4 ? offset_211 : _GEN_6392; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7429 = _T_4 ? offset_212 : _GEN_6393; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7430 = _T_4 ? offset_213 : _GEN_6394; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7431 = _T_4 ? offset_214 : _GEN_6395; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7432 = _T_4 ? offset_215 : _GEN_6396; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7433 = _T_4 ? offset_216 : _GEN_6397; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7434 = _T_4 ? offset_217 : _GEN_6398; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7435 = _T_4 ? offset_218 : _GEN_6399; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7436 = _T_4 ? offset_219 : _GEN_6400; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7437 = _T_4 ? offset_220 : _GEN_6401; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7438 = _T_4 ? offset_221 : _GEN_6402; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7439 = _T_4 ? offset_222 : _GEN_6403; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7440 = _T_4 ? offset_223 : _GEN_6404; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7441 = _T_4 ? offset_224 : _GEN_6405; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7442 = _T_4 ? offset_225 : _GEN_6406; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7443 = _T_4 ? offset_226 : _GEN_6407; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7444 = _T_4 ? offset_227 : _GEN_6408; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7445 = _T_4 ? offset_228 : _GEN_6409; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7446 = _T_4 ? offset_229 : _GEN_6410; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7447 = _T_4 ? offset_230 : _GEN_6411; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7448 = _T_4 ? offset_231 : _GEN_6412; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7449 = _T_4 ? offset_232 : _GEN_6413; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7450 = _T_4 ? offset_233 : _GEN_6414; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7451 = _T_4 ? offset_234 : _GEN_6415; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7452 = _T_4 ? offset_235 : _GEN_6416; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7453 = _T_4 ? offset_236 : _GEN_6417; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7454 = _T_4 ? offset_237 : _GEN_6418; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7455 = _T_4 ? offset_238 : _GEN_6419; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7456 = _T_4 ? offset_239 : _GEN_6420; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7457 = _T_4 ? offset_240 : _GEN_6421; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7458 = _T_4 ? offset_241 : _GEN_6422; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7459 = _T_4 ? offset_242 : _GEN_6423; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7460 = _T_4 ? offset_243 : _GEN_6424; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7461 = _T_4 ? offset_244 : _GEN_6425; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7462 = _T_4 ? offset_245 : _GEN_6426; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7463 = _T_4 ? offset_246 : _GEN_6427; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7464 = _T_4 ? offset_247 : _GEN_6428; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7465 = _T_4 ? offset_248 : _GEN_6429; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7466 = _T_4 ? offset_249 : _GEN_6430; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7467 = _T_4 ? offset_250 : _GEN_6431; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7468 = _T_4 ? offset_251 : _GEN_6432; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7469 = _T_4 ? offset_252 : _GEN_6433; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7470 = _T_4 ? offset_253 : _GEN_6434; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7471 = _T_4 ? offset_254 : _GEN_6435; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [3:0] _GEN_7472 = _T_4 ? offset_255 : _GEN_6436; // @[Conditional.scala 39:67 Dcache.scala 19:24]
  wire [31:0] _GEN_7473 = _T_3 ? _data_addr_T : _GEN_6438; // @[Conditional.scala 39:67 Dcache.scala 153:21]
  wire [127:0] _GEN_7474 = _T_3 ? cache_data_out : 128'h0; // @[Conditional.scala 39:67 Dcache.scala 154:21]
  wire [7:0] _GEN_7475 = _T_3 ? 8'hff : 8'h0; // @[Conditional.scala 39:67 Dcache.scala 155:21]
  wire  _GEN_7477 = _T_3 ? _GEN_3336 : _GEN_6442; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_9538 = _T_1 ? 32'h0 : _GEN_7473; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_9539 = _T_1 ? 128'h0 : _GEN_7474; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_9540 = _T_1 ? 8'h0 : _GEN_7475; // @[Conditional.scala 39:67]
  wire  _GEN_9542 = _T_1 ? 1'h0 : _GEN_7477; // @[Conditional.scala 39:67]
  wire  _GEN_9543 = _T_1 ? 1'h0 : _T_3 & _GEN_3336; // @[Conditional.scala 39:67]
  S011HD1P_X32Y2D128_BW req ( // @[Dcache.scala 217:19]
    .Q(req_Q),
    .CLK(req_CLK),
    .CEN(req_CEN),
    .WEN(req_WEN),
    .BWEN(req_BWEN),
    .A(req_A),
    .D(req_D)
  );
  assign io_dmem_data_ready = data_ready; // @[Dcache.scala 214:19]
  assign io_dmem_data_read = 2'h3 == io_dmem_data_size ? valid_rdata : {{31'd0}, _data_read_T_42}; // @[Mux.scala 80:57]
  assign io_out_data_valid = _T ? 1'h0 : _GEN_9542; // @[Conditional.scala 40:58]
  assign io_out_data_req = _T ? 1'h0 : _GEN_9543; // @[Conditional.scala 40:58]
  assign io_out_data_addr = _T ? 32'h0 : _GEN_9538; // @[Conditional.scala 40:58]
  assign io_out_data_strb = _T ? 8'h0 : _GEN_9540; // @[Conditional.scala 40:58]
  assign io_out_data_write = _T ? 128'h0 : _GEN_9539; // @[Conditional.scala 40:58]
  assign req_CLK = clock; // @[Dcache.scala 218:17]
  assign req_CEN = 1'h1; // @[Dcache.scala 219:17]
  assign req_WEN = cache_wen; // @[Dcache.scala 220:17]
  assign req_BWEN = cache_strb; // @[Dcache.scala 221:17]
  assign req_A = io_dmem_data_addr[11:4]; // @[Dcache.scala 29:30]
  assign req_D = cache_wdata; // @[Dcache.scala 223:17]
  always @(posedge clock) begin
    if (reset) begin // @[Dcache.scala 16:24]
      tag_0 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_0 <= _GEN_1025;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_0 <= _GEN_6705;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_1 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_1 <= _GEN_1026;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_1 <= _GEN_6706;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_2 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_2 <= _GEN_1027;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_2 <= _GEN_6707;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_3 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_3 <= _GEN_1028;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_3 <= _GEN_6708;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_4 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_4 <= _GEN_1029;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_4 <= _GEN_6709;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_5 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_5 <= _GEN_1030;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_5 <= _GEN_6710;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_6 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_6 <= _GEN_1031;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_6 <= _GEN_6711;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_7 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_7 <= _GEN_1032;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_7 <= _GEN_6712;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_8 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_8 <= _GEN_1033;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_8 <= _GEN_6713;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_9 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_9 <= _GEN_1034;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_9 <= _GEN_6714;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_10 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_10 <= _GEN_1035;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_10 <= _GEN_6715;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_11 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_11 <= _GEN_1036;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_11 <= _GEN_6716;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_12 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_12 <= _GEN_1037;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_12 <= _GEN_6717;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_13 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_13 <= _GEN_1038;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_13 <= _GEN_6718;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_14 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_14 <= _GEN_1039;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_14 <= _GEN_6719;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_15 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_15 <= _GEN_1040;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_15 <= _GEN_6720;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_16 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_16 <= _GEN_1041;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_16 <= _GEN_6721;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_17 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_17 <= _GEN_1042;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_17 <= _GEN_6722;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_18 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_18 <= _GEN_1043;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_18 <= _GEN_6723;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_19 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_19 <= _GEN_1044;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_19 <= _GEN_6724;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_20 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_20 <= _GEN_1045;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_20 <= _GEN_6725;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_21 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_21 <= _GEN_1046;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_21 <= _GEN_6726;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_22 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_22 <= _GEN_1047;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_22 <= _GEN_6727;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_23 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_23 <= _GEN_1048;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_23 <= _GEN_6728;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_24 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_24 <= _GEN_1049;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_24 <= _GEN_6729;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_25 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_25 <= _GEN_1050;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_25 <= _GEN_6730;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_26 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_26 <= _GEN_1051;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_26 <= _GEN_6731;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_27 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_27 <= _GEN_1052;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_27 <= _GEN_6732;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_28 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_28 <= _GEN_1053;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_28 <= _GEN_6733;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_29 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_29 <= _GEN_1054;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_29 <= _GEN_6734;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_30 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_30 <= _GEN_1055;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_30 <= _GEN_6735;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_31 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_31 <= _GEN_1056;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_31 <= _GEN_6736;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_32 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_32 <= _GEN_1057;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_32 <= _GEN_6737;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_33 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_33 <= _GEN_1058;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_33 <= _GEN_6738;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_34 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_34 <= _GEN_1059;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_34 <= _GEN_6739;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_35 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_35 <= _GEN_1060;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_35 <= _GEN_6740;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_36 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_36 <= _GEN_1061;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_36 <= _GEN_6741;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_37 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_37 <= _GEN_1062;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_37 <= _GEN_6742;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_38 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_38 <= _GEN_1063;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_38 <= _GEN_6743;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_39 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_39 <= _GEN_1064;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_39 <= _GEN_6744;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_40 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_40 <= _GEN_1065;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_40 <= _GEN_6745;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_41 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_41 <= _GEN_1066;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_41 <= _GEN_6746;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_42 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_42 <= _GEN_1067;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_42 <= _GEN_6747;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_43 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_43 <= _GEN_1068;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_43 <= _GEN_6748;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_44 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_44 <= _GEN_1069;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_44 <= _GEN_6749;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_45 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_45 <= _GEN_1070;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_45 <= _GEN_6750;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_46 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_46 <= _GEN_1071;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_46 <= _GEN_6751;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_47 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_47 <= _GEN_1072;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_47 <= _GEN_6752;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_48 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_48 <= _GEN_1073;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_48 <= _GEN_6753;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_49 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_49 <= _GEN_1074;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_49 <= _GEN_6754;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_50 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_50 <= _GEN_1075;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_50 <= _GEN_6755;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_51 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_51 <= _GEN_1076;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_51 <= _GEN_6756;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_52 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_52 <= _GEN_1077;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_52 <= _GEN_6757;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_53 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_53 <= _GEN_1078;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_53 <= _GEN_6758;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_54 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_54 <= _GEN_1079;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_54 <= _GEN_6759;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_55 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_55 <= _GEN_1080;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_55 <= _GEN_6760;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_56 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_56 <= _GEN_1081;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_56 <= _GEN_6761;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_57 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_57 <= _GEN_1082;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_57 <= _GEN_6762;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_58 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_58 <= _GEN_1083;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_58 <= _GEN_6763;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_59 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_59 <= _GEN_1084;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_59 <= _GEN_6764;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_60 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_60 <= _GEN_1085;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_60 <= _GEN_6765;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_61 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_61 <= _GEN_1086;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_61 <= _GEN_6766;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_62 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_62 <= _GEN_1087;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_62 <= _GEN_6767;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_63 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_63 <= _GEN_1088;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_63 <= _GEN_6768;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_64 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_64 <= _GEN_1089;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_64 <= _GEN_6769;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_65 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_65 <= _GEN_1090;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_65 <= _GEN_6770;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_66 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_66 <= _GEN_1091;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_66 <= _GEN_6771;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_67 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_67 <= _GEN_1092;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_67 <= _GEN_6772;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_68 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_68 <= _GEN_1093;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_68 <= _GEN_6773;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_69 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_69 <= _GEN_1094;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_69 <= _GEN_6774;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_70 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_70 <= _GEN_1095;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_70 <= _GEN_6775;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_71 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_71 <= _GEN_1096;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_71 <= _GEN_6776;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_72 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_72 <= _GEN_1097;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_72 <= _GEN_6777;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_73 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_73 <= _GEN_1098;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_73 <= _GEN_6778;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_74 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_74 <= _GEN_1099;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_74 <= _GEN_6779;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_75 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_75 <= _GEN_1100;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_75 <= _GEN_6780;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_76 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_76 <= _GEN_1101;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_76 <= _GEN_6781;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_77 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_77 <= _GEN_1102;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_77 <= _GEN_6782;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_78 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_78 <= _GEN_1103;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_78 <= _GEN_6783;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_79 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_79 <= _GEN_1104;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_79 <= _GEN_6784;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_80 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_80 <= _GEN_1105;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_80 <= _GEN_6785;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_81 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_81 <= _GEN_1106;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_81 <= _GEN_6786;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_82 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_82 <= _GEN_1107;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_82 <= _GEN_6787;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_83 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_83 <= _GEN_1108;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_83 <= _GEN_6788;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_84 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_84 <= _GEN_1109;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_84 <= _GEN_6789;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_85 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_85 <= _GEN_1110;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_85 <= _GEN_6790;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_86 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_86 <= _GEN_1111;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_86 <= _GEN_6791;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_87 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_87 <= _GEN_1112;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_87 <= _GEN_6792;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_88 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_88 <= _GEN_1113;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_88 <= _GEN_6793;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_89 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_89 <= _GEN_1114;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_89 <= _GEN_6794;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_90 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_90 <= _GEN_1115;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_90 <= _GEN_6795;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_91 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_91 <= _GEN_1116;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_91 <= _GEN_6796;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_92 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_92 <= _GEN_1117;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_92 <= _GEN_6797;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_93 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_93 <= _GEN_1118;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_93 <= _GEN_6798;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_94 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_94 <= _GEN_1119;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_94 <= _GEN_6799;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_95 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_95 <= _GEN_1120;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_95 <= _GEN_6800;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_96 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_96 <= _GEN_1121;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_96 <= _GEN_6801;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_97 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_97 <= _GEN_1122;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_97 <= _GEN_6802;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_98 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_98 <= _GEN_1123;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_98 <= _GEN_6803;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_99 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_99 <= _GEN_1124;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_99 <= _GEN_6804;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_100 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_100 <= _GEN_1125;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_100 <= _GEN_6805;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_101 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_101 <= _GEN_1126;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_101 <= _GEN_6806;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_102 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_102 <= _GEN_1127;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_102 <= _GEN_6807;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_103 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_103 <= _GEN_1128;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_103 <= _GEN_6808;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_104 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_104 <= _GEN_1129;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_104 <= _GEN_6809;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_105 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_105 <= _GEN_1130;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_105 <= _GEN_6810;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_106 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_106 <= _GEN_1131;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_106 <= _GEN_6811;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_107 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_107 <= _GEN_1132;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_107 <= _GEN_6812;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_108 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_108 <= _GEN_1133;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_108 <= _GEN_6813;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_109 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_109 <= _GEN_1134;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_109 <= _GEN_6814;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_110 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_110 <= _GEN_1135;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_110 <= _GEN_6815;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_111 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_111 <= _GEN_1136;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_111 <= _GEN_6816;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_112 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_112 <= _GEN_1137;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_112 <= _GEN_6817;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_113 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_113 <= _GEN_1138;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_113 <= _GEN_6818;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_114 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_114 <= _GEN_1139;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_114 <= _GEN_6819;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_115 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_115 <= _GEN_1140;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_115 <= _GEN_6820;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_116 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_116 <= _GEN_1141;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_116 <= _GEN_6821;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_117 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_117 <= _GEN_1142;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_117 <= _GEN_6822;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_118 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_118 <= _GEN_1143;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_118 <= _GEN_6823;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_119 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_119 <= _GEN_1144;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_119 <= _GEN_6824;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_120 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_120 <= _GEN_1145;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_120 <= _GEN_6825;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_121 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_121 <= _GEN_1146;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_121 <= _GEN_6826;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_122 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_122 <= _GEN_1147;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_122 <= _GEN_6827;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_123 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_123 <= _GEN_1148;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_123 <= _GEN_6828;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_124 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_124 <= _GEN_1149;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_124 <= _GEN_6829;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_125 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_125 <= _GEN_1150;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_125 <= _GEN_6830;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_126 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_126 <= _GEN_1151;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_126 <= _GEN_6831;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_127 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_127 <= _GEN_1152;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_127 <= _GEN_6832;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_128 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_128 <= _GEN_1153;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_128 <= _GEN_6833;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_129 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_129 <= _GEN_1154;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_129 <= _GEN_6834;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_130 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_130 <= _GEN_1155;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_130 <= _GEN_6835;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_131 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_131 <= _GEN_1156;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_131 <= _GEN_6836;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_132 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_132 <= _GEN_1157;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_132 <= _GEN_6837;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_133 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_133 <= _GEN_1158;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_133 <= _GEN_6838;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_134 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_134 <= _GEN_1159;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_134 <= _GEN_6839;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_135 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_135 <= _GEN_1160;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_135 <= _GEN_6840;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_136 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_136 <= _GEN_1161;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_136 <= _GEN_6841;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_137 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_137 <= _GEN_1162;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_137 <= _GEN_6842;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_138 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_138 <= _GEN_1163;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_138 <= _GEN_6843;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_139 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_139 <= _GEN_1164;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_139 <= _GEN_6844;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_140 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_140 <= _GEN_1165;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_140 <= _GEN_6845;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_141 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_141 <= _GEN_1166;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_141 <= _GEN_6846;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_142 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_142 <= _GEN_1167;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_142 <= _GEN_6847;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_143 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_143 <= _GEN_1168;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_143 <= _GEN_6848;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_144 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_144 <= _GEN_1169;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_144 <= _GEN_6849;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_145 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_145 <= _GEN_1170;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_145 <= _GEN_6850;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_146 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_146 <= _GEN_1171;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_146 <= _GEN_6851;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_147 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_147 <= _GEN_1172;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_147 <= _GEN_6852;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_148 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_148 <= _GEN_1173;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_148 <= _GEN_6853;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_149 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_149 <= _GEN_1174;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_149 <= _GEN_6854;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_150 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_150 <= _GEN_1175;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_150 <= _GEN_6855;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_151 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_151 <= _GEN_1176;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_151 <= _GEN_6856;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_152 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_152 <= _GEN_1177;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_152 <= _GEN_6857;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_153 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_153 <= _GEN_1178;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_153 <= _GEN_6858;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_154 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_154 <= _GEN_1179;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_154 <= _GEN_6859;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_155 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_155 <= _GEN_1180;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_155 <= _GEN_6860;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_156 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_156 <= _GEN_1181;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_156 <= _GEN_6861;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_157 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_157 <= _GEN_1182;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_157 <= _GEN_6862;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_158 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_158 <= _GEN_1183;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_158 <= _GEN_6863;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_159 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_159 <= _GEN_1184;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_159 <= _GEN_6864;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_160 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_160 <= _GEN_1185;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_160 <= _GEN_6865;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_161 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_161 <= _GEN_1186;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_161 <= _GEN_6866;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_162 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_162 <= _GEN_1187;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_162 <= _GEN_6867;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_163 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_163 <= _GEN_1188;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_163 <= _GEN_6868;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_164 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_164 <= _GEN_1189;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_164 <= _GEN_6869;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_165 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_165 <= _GEN_1190;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_165 <= _GEN_6870;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_166 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_166 <= _GEN_1191;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_166 <= _GEN_6871;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_167 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_167 <= _GEN_1192;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_167 <= _GEN_6872;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_168 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_168 <= _GEN_1193;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_168 <= _GEN_6873;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_169 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_169 <= _GEN_1194;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_169 <= _GEN_6874;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_170 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_170 <= _GEN_1195;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_170 <= _GEN_6875;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_171 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_171 <= _GEN_1196;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_171 <= _GEN_6876;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_172 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_172 <= _GEN_1197;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_172 <= _GEN_6877;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_173 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_173 <= _GEN_1198;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_173 <= _GEN_6878;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_174 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_174 <= _GEN_1199;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_174 <= _GEN_6879;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_175 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_175 <= _GEN_1200;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_175 <= _GEN_6880;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_176 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_176 <= _GEN_1201;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_176 <= _GEN_6881;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_177 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_177 <= _GEN_1202;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_177 <= _GEN_6882;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_178 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_178 <= _GEN_1203;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_178 <= _GEN_6883;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_179 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_179 <= _GEN_1204;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_179 <= _GEN_6884;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_180 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_180 <= _GEN_1205;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_180 <= _GEN_6885;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_181 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_181 <= _GEN_1206;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_181 <= _GEN_6886;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_182 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_182 <= _GEN_1207;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_182 <= _GEN_6887;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_183 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_183 <= _GEN_1208;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_183 <= _GEN_6888;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_184 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_184 <= _GEN_1209;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_184 <= _GEN_6889;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_185 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_185 <= _GEN_1210;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_185 <= _GEN_6890;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_186 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_186 <= _GEN_1211;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_186 <= _GEN_6891;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_187 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_187 <= _GEN_1212;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_187 <= _GEN_6892;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_188 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_188 <= _GEN_1213;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_188 <= _GEN_6893;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_189 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_189 <= _GEN_1214;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_189 <= _GEN_6894;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_190 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_190 <= _GEN_1215;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_190 <= _GEN_6895;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_191 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_191 <= _GEN_1216;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_191 <= _GEN_6896;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_192 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_192 <= _GEN_1217;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_192 <= _GEN_6897;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_193 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_193 <= _GEN_1218;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_193 <= _GEN_6898;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_194 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_194 <= _GEN_1219;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_194 <= _GEN_6899;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_195 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_195 <= _GEN_1220;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_195 <= _GEN_6900;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_196 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_196 <= _GEN_1221;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_196 <= _GEN_6901;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_197 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_197 <= _GEN_1222;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_197 <= _GEN_6902;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_198 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_198 <= _GEN_1223;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_198 <= _GEN_6903;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_199 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_199 <= _GEN_1224;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_199 <= _GEN_6904;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_200 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_200 <= _GEN_1225;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_200 <= _GEN_6905;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_201 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_201 <= _GEN_1226;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_201 <= _GEN_6906;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_202 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_202 <= _GEN_1227;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_202 <= _GEN_6907;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_203 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_203 <= _GEN_1228;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_203 <= _GEN_6908;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_204 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_204 <= _GEN_1229;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_204 <= _GEN_6909;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_205 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_205 <= _GEN_1230;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_205 <= _GEN_6910;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_206 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_206 <= _GEN_1231;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_206 <= _GEN_6911;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_207 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_207 <= _GEN_1232;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_207 <= _GEN_6912;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_208 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_208 <= _GEN_1233;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_208 <= _GEN_6913;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_209 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_209 <= _GEN_1234;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_209 <= _GEN_6914;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_210 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_210 <= _GEN_1235;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_210 <= _GEN_6915;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_211 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_211 <= _GEN_1236;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_211 <= _GEN_6916;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_212 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_212 <= _GEN_1237;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_212 <= _GEN_6917;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_213 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_213 <= _GEN_1238;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_213 <= _GEN_6918;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_214 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_214 <= _GEN_1239;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_214 <= _GEN_6919;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_215 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_215 <= _GEN_1240;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_215 <= _GEN_6920;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_216 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_216 <= _GEN_1241;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_216 <= _GEN_6921;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_217 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_217 <= _GEN_1242;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_217 <= _GEN_6922;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_218 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_218 <= _GEN_1243;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_218 <= _GEN_6923;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_219 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_219 <= _GEN_1244;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_219 <= _GEN_6924;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_220 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_220 <= _GEN_1245;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_220 <= _GEN_6925;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_221 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_221 <= _GEN_1246;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_221 <= _GEN_6926;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_222 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_222 <= _GEN_1247;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_222 <= _GEN_6927;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_223 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_223 <= _GEN_1248;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_223 <= _GEN_6928;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_224 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_224 <= _GEN_1249;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_224 <= _GEN_6929;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_225 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_225 <= _GEN_1250;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_225 <= _GEN_6930;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_226 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_226 <= _GEN_1251;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_226 <= _GEN_6931;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_227 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_227 <= _GEN_1252;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_227 <= _GEN_6932;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_228 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_228 <= _GEN_1253;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_228 <= _GEN_6933;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_229 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_229 <= _GEN_1254;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_229 <= _GEN_6934;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_230 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_230 <= _GEN_1255;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_230 <= _GEN_6935;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_231 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_231 <= _GEN_1256;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_231 <= _GEN_6936;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_232 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_232 <= _GEN_1257;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_232 <= _GEN_6937;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_233 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_233 <= _GEN_1258;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_233 <= _GEN_6938;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_234 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_234 <= _GEN_1259;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_234 <= _GEN_6939;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_235 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_235 <= _GEN_1260;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_235 <= _GEN_6940;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_236 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_236 <= _GEN_1261;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_236 <= _GEN_6941;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_237 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_237 <= _GEN_1262;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_237 <= _GEN_6942;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_238 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_238 <= _GEN_1263;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_238 <= _GEN_6943;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_239 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_239 <= _GEN_1264;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_239 <= _GEN_6944;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_240 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_240 <= _GEN_1265;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_240 <= _GEN_6945;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_241 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_241 <= _GEN_1266;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_241 <= _GEN_6946;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_242 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_242 <= _GEN_1267;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_242 <= _GEN_6947;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_243 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_243 <= _GEN_1268;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_243 <= _GEN_6948;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_244 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_244 <= _GEN_1269;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_244 <= _GEN_6949;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_245 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_245 <= _GEN_1270;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_245 <= _GEN_6950;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_246 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_246 <= _GEN_1271;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_246 <= _GEN_6951;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_247 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_247 <= _GEN_1272;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_247 <= _GEN_6952;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_248 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_248 <= _GEN_1273;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_248 <= _GEN_6953;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_249 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_249 <= _GEN_1274;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_249 <= _GEN_6954;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_250 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_250 <= _GEN_1275;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_250 <= _GEN_6955;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_251 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_251 <= _GEN_1276;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_251 <= _GEN_6956;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_252 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_252 <= _GEN_1277;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_252 <= _GEN_6957;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_253 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_253 <= _GEN_1278;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_253 <= _GEN_6958;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_254 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_254 <= _GEN_1279;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_254 <= _GEN_6959;
      end
    end
    if (reset) begin // @[Dcache.scala 16:24]
      tag_255 <= 20'h0; // @[Dcache.scala 16:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          tag_255 <= _GEN_1280;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        tag_255 <= _GEN_6960;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_0 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_0 <= _GEN_769;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_0 <= _GEN_6449;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_1 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_1 <= _GEN_770;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_1 <= _GEN_6450;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_2 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_2 <= _GEN_771;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_2 <= _GEN_6451;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_3 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_3 <= _GEN_772;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_3 <= _GEN_6452;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_4 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_4 <= _GEN_773;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_4 <= _GEN_6453;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_5 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_5 <= _GEN_774;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_5 <= _GEN_6454;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_6 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_6 <= _GEN_775;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_6 <= _GEN_6455;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_7 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_7 <= _GEN_776;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_7 <= _GEN_6456;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_8 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_8 <= _GEN_777;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_8 <= _GEN_6457;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_9 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_9 <= _GEN_778;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_9 <= _GEN_6458;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_10 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_10 <= _GEN_779;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_10 <= _GEN_6459;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_11 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_11 <= _GEN_780;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_11 <= _GEN_6460;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_12 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_12 <= _GEN_781;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_12 <= _GEN_6461;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_13 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_13 <= _GEN_782;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_13 <= _GEN_6462;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_14 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_14 <= _GEN_783;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_14 <= _GEN_6463;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_15 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_15 <= _GEN_784;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_15 <= _GEN_6464;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_16 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_16 <= _GEN_785;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_16 <= _GEN_6465;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_17 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_17 <= _GEN_786;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_17 <= _GEN_6466;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_18 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_18 <= _GEN_787;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_18 <= _GEN_6467;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_19 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_19 <= _GEN_788;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_19 <= _GEN_6468;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_20 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_20 <= _GEN_789;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_20 <= _GEN_6469;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_21 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_21 <= _GEN_790;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_21 <= _GEN_6470;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_22 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_22 <= _GEN_791;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_22 <= _GEN_6471;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_23 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_23 <= _GEN_792;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_23 <= _GEN_6472;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_24 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_24 <= _GEN_793;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_24 <= _GEN_6473;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_25 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_25 <= _GEN_794;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_25 <= _GEN_6474;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_26 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_26 <= _GEN_795;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_26 <= _GEN_6475;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_27 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_27 <= _GEN_796;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_27 <= _GEN_6476;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_28 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_28 <= _GEN_797;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_28 <= _GEN_6477;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_29 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_29 <= _GEN_798;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_29 <= _GEN_6478;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_30 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_30 <= _GEN_799;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_30 <= _GEN_6479;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_31 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_31 <= _GEN_800;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_31 <= _GEN_6480;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_32 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_32 <= _GEN_801;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_32 <= _GEN_6481;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_33 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_33 <= _GEN_802;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_33 <= _GEN_6482;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_34 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_34 <= _GEN_803;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_34 <= _GEN_6483;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_35 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_35 <= _GEN_804;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_35 <= _GEN_6484;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_36 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_36 <= _GEN_805;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_36 <= _GEN_6485;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_37 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_37 <= _GEN_806;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_37 <= _GEN_6486;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_38 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_38 <= _GEN_807;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_38 <= _GEN_6487;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_39 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_39 <= _GEN_808;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_39 <= _GEN_6488;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_40 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_40 <= _GEN_809;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_40 <= _GEN_6489;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_41 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_41 <= _GEN_810;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_41 <= _GEN_6490;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_42 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_42 <= _GEN_811;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_42 <= _GEN_6491;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_43 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_43 <= _GEN_812;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_43 <= _GEN_6492;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_44 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_44 <= _GEN_813;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_44 <= _GEN_6493;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_45 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_45 <= _GEN_814;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_45 <= _GEN_6494;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_46 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_46 <= _GEN_815;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_46 <= _GEN_6495;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_47 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_47 <= _GEN_816;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_47 <= _GEN_6496;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_48 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_48 <= _GEN_817;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_48 <= _GEN_6497;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_49 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_49 <= _GEN_818;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_49 <= _GEN_6498;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_50 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_50 <= _GEN_819;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_50 <= _GEN_6499;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_51 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_51 <= _GEN_820;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_51 <= _GEN_6500;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_52 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_52 <= _GEN_821;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_52 <= _GEN_6501;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_53 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_53 <= _GEN_822;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_53 <= _GEN_6502;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_54 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_54 <= _GEN_823;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_54 <= _GEN_6503;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_55 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_55 <= _GEN_824;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_55 <= _GEN_6504;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_56 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_56 <= _GEN_825;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_56 <= _GEN_6505;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_57 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_57 <= _GEN_826;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_57 <= _GEN_6506;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_58 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_58 <= _GEN_827;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_58 <= _GEN_6507;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_59 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_59 <= _GEN_828;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_59 <= _GEN_6508;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_60 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_60 <= _GEN_829;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_60 <= _GEN_6509;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_61 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_61 <= _GEN_830;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_61 <= _GEN_6510;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_62 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_62 <= _GEN_831;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_62 <= _GEN_6511;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_63 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_63 <= _GEN_832;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_63 <= _GEN_6512;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_64 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_64 <= _GEN_833;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_64 <= _GEN_6513;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_65 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_65 <= _GEN_834;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_65 <= _GEN_6514;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_66 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_66 <= _GEN_835;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_66 <= _GEN_6515;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_67 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_67 <= _GEN_836;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_67 <= _GEN_6516;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_68 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_68 <= _GEN_837;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_68 <= _GEN_6517;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_69 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_69 <= _GEN_838;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_69 <= _GEN_6518;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_70 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_70 <= _GEN_839;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_70 <= _GEN_6519;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_71 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_71 <= _GEN_840;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_71 <= _GEN_6520;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_72 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_72 <= _GEN_841;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_72 <= _GEN_6521;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_73 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_73 <= _GEN_842;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_73 <= _GEN_6522;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_74 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_74 <= _GEN_843;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_74 <= _GEN_6523;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_75 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_75 <= _GEN_844;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_75 <= _GEN_6524;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_76 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_76 <= _GEN_845;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_76 <= _GEN_6525;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_77 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_77 <= _GEN_846;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_77 <= _GEN_6526;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_78 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_78 <= _GEN_847;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_78 <= _GEN_6527;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_79 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_79 <= _GEN_848;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_79 <= _GEN_6528;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_80 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_80 <= _GEN_849;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_80 <= _GEN_6529;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_81 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_81 <= _GEN_850;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_81 <= _GEN_6530;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_82 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_82 <= _GEN_851;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_82 <= _GEN_6531;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_83 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_83 <= _GEN_852;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_83 <= _GEN_6532;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_84 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_84 <= _GEN_853;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_84 <= _GEN_6533;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_85 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_85 <= _GEN_854;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_85 <= _GEN_6534;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_86 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_86 <= _GEN_855;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_86 <= _GEN_6535;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_87 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_87 <= _GEN_856;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_87 <= _GEN_6536;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_88 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_88 <= _GEN_857;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_88 <= _GEN_6537;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_89 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_89 <= _GEN_858;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_89 <= _GEN_6538;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_90 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_90 <= _GEN_859;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_90 <= _GEN_6539;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_91 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_91 <= _GEN_860;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_91 <= _GEN_6540;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_92 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_92 <= _GEN_861;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_92 <= _GEN_6541;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_93 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_93 <= _GEN_862;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_93 <= _GEN_6542;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_94 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_94 <= _GEN_863;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_94 <= _GEN_6543;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_95 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_95 <= _GEN_864;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_95 <= _GEN_6544;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_96 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_96 <= _GEN_865;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_96 <= _GEN_6545;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_97 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_97 <= _GEN_866;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_97 <= _GEN_6546;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_98 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_98 <= _GEN_867;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_98 <= _GEN_6547;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_99 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_99 <= _GEN_868;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_99 <= _GEN_6548;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_100 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_100 <= _GEN_869;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_100 <= _GEN_6549;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_101 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_101 <= _GEN_870;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_101 <= _GEN_6550;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_102 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_102 <= _GEN_871;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_102 <= _GEN_6551;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_103 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_103 <= _GEN_872;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_103 <= _GEN_6552;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_104 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_104 <= _GEN_873;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_104 <= _GEN_6553;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_105 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_105 <= _GEN_874;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_105 <= _GEN_6554;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_106 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_106 <= _GEN_875;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_106 <= _GEN_6555;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_107 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_107 <= _GEN_876;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_107 <= _GEN_6556;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_108 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_108 <= _GEN_877;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_108 <= _GEN_6557;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_109 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_109 <= _GEN_878;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_109 <= _GEN_6558;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_110 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_110 <= _GEN_879;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_110 <= _GEN_6559;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_111 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_111 <= _GEN_880;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_111 <= _GEN_6560;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_112 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_112 <= _GEN_881;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_112 <= _GEN_6561;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_113 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_113 <= _GEN_882;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_113 <= _GEN_6562;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_114 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_114 <= _GEN_883;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_114 <= _GEN_6563;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_115 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_115 <= _GEN_884;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_115 <= _GEN_6564;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_116 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_116 <= _GEN_885;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_116 <= _GEN_6565;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_117 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_117 <= _GEN_886;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_117 <= _GEN_6566;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_118 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_118 <= _GEN_887;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_118 <= _GEN_6567;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_119 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_119 <= _GEN_888;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_119 <= _GEN_6568;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_120 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_120 <= _GEN_889;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_120 <= _GEN_6569;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_121 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_121 <= _GEN_890;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_121 <= _GEN_6570;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_122 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_122 <= _GEN_891;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_122 <= _GEN_6571;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_123 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_123 <= _GEN_892;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_123 <= _GEN_6572;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_124 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_124 <= _GEN_893;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_124 <= _GEN_6573;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_125 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_125 <= _GEN_894;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_125 <= _GEN_6574;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_126 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_126 <= _GEN_895;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_126 <= _GEN_6575;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_127 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_127 <= _GEN_896;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_127 <= _GEN_6576;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_128 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_128 <= _GEN_897;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_128 <= _GEN_6577;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_129 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_129 <= _GEN_898;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_129 <= _GEN_6578;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_130 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_130 <= _GEN_899;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_130 <= _GEN_6579;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_131 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_131 <= _GEN_900;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_131 <= _GEN_6580;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_132 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_132 <= _GEN_901;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_132 <= _GEN_6581;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_133 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_133 <= _GEN_902;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_133 <= _GEN_6582;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_134 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_134 <= _GEN_903;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_134 <= _GEN_6583;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_135 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_135 <= _GEN_904;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_135 <= _GEN_6584;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_136 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_136 <= _GEN_905;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_136 <= _GEN_6585;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_137 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_137 <= _GEN_906;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_137 <= _GEN_6586;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_138 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_138 <= _GEN_907;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_138 <= _GEN_6587;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_139 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_139 <= _GEN_908;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_139 <= _GEN_6588;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_140 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_140 <= _GEN_909;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_140 <= _GEN_6589;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_141 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_141 <= _GEN_910;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_141 <= _GEN_6590;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_142 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_142 <= _GEN_911;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_142 <= _GEN_6591;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_143 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_143 <= _GEN_912;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_143 <= _GEN_6592;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_144 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_144 <= _GEN_913;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_144 <= _GEN_6593;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_145 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_145 <= _GEN_914;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_145 <= _GEN_6594;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_146 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_146 <= _GEN_915;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_146 <= _GEN_6595;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_147 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_147 <= _GEN_916;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_147 <= _GEN_6596;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_148 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_148 <= _GEN_917;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_148 <= _GEN_6597;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_149 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_149 <= _GEN_918;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_149 <= _GEN_6598;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_150 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_150 <= _GEN_919;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_150 <= _GEN_6599;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_151 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_151 <= _GEN_920;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_151 <= _GEN_6600;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_152 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_152 <= _GEN_921;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_152 <= _GEN_6601;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_153 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_153 <= _GEN_922;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_153 <= _GEN_6602;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_154 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_154 <= _GEN_923;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_154 <= _GEN_6603;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_155 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_155 <= _GEN_924;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_155 <= _GEN_6604;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_156 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_156 <= _GEN_925;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_156 <= _GEN_6605;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_157 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_157 <= _GEN_926;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_157 <= _GEN_6606;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_158 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_158 <= _GEN_927;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_158 <= _GEN_6607;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_159 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_159 <= _GEN_928;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_159 <= _GEN_6608;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_160 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_160 <= _GEN_929;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_160 <= _GEN_6609;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_161 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_161 <= _GEN_930;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_161 <= _GEN_6610;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_162 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_162 <= _GEN_931;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_162 <= _GEN_6611;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_163 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_163 <= _GEN_932;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_163 <= _GEN_6612;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_164 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_164 <= _GEN_933;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_164 <= _GEN_6613;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_165 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_165 <= _GEN_934;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_165 <= _GEN_6614;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_166 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_166 <= _GEN_935;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_166 <= _GEN_6615;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_167 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_167 <= _GEN_936;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_167 <= _GEN_6616;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_168 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_168 <= _GEN_937;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_168 <= _GEN_6617;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_169 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_169 <= _GEN_938;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_169 <= _GEN_6618;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_170 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_170 <= _GEN_939;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_170 <= _GEN_6619;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_171 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_171 <= _GEN_940;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_171 <= _GEN_6620;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_172 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_172 <= _GEN_941;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_172 <= _GEN_6621;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_173 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_173 <= _GEN_942;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_173 <= _GEN_6622;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_174 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_174 <= _GEN_943;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_174 <= _GEN_6623;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_175 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_175 <= _GEN_944;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_175 <= _GEN_6624;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_176 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_176 <= _GEN_945;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_176 <= _GEN_6625;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_177 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_177 <= _GEN_946;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_177 <= _GEN_6626;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_178 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_178 <= _GEN_947;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_178 <= _GEN_6627;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_179 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_179 <= _GEN_948;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_179 <= _GEN_6628;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_180 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_180 <= _GEN_949;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_180 <= _GEN_6629;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_181 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_181 <= _GEN_950;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_181 <= _GEN_6630;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_182 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_182 <= _GEN_951;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_182 <= _GEN_6631;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_183 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_183 <= _GEN_952;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_183 <= _GEN_6632;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_184 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_184 <= _GEN_953;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_184 <= _GEN_6633;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_185 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_185 <= _GEN_954;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_185 <= _GEN_6634;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_186 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_186 <= _GEN_955;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_186 <= _GEN_6635;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_187 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_187 <= _GEN_956;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_187 <= _GEN_6636;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_188 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_188 <= _GEN_957;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_188 <= _GEN_6637;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_189 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_189 <= _GEN_958;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_189 <= _GEN_6638;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_190 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_190 <= _GEN_959;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_190 <= _GEN_6639;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_191 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_191 <= _GEN_960;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_191 <= _GEN_6640;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_192 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_192 <= _GEN_961;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_192 <= _GEN_6641;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_193 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_193 <= _GEN_962;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_193 <= _GEN_6642;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_194 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_194 <= _GEN_963;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_194 <= _GEN_6643;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_195 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_195 <= _GEN_964;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_195 <= _GEN_6644;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_196 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_196 <= _GEN_965;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_196 <= _GEN_6645;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_197 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_197 <= _GEN_966;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_197 <= _GEN_6646;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_198 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_198 <= _GEN_967;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_198 <= _GEN_6647;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_199 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_199 <= _GEN_968;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_199 <= _GEN_6648;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_200 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_200 <= _GEN_969;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_200 <= _GEN_6649;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_201 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_201 <= _GEN_970;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_201 <= _GEN_6650;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_202 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_202 <= _GEN_971;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_202 <= _GEN_6651;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_203 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_203 <= _GEN_972;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_203 <= _GEN_6652;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_204 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_204 <= _GEN_973;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_204 <= _GEN_6653;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_205 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_205 <= _GEN_974;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_205 <= _GEN_6654;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_206 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_206 <= _GEN_975;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_206 <= _GEN_6655;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_207 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_207 <= _GEN_976;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_207 <= _GEN_6656;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_208 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_208 <= _GEN_977;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_208 <= _GEN_6657;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_209 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_209 <= _GEN_978;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_209 <= _GEN_6658;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_210 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_210 <= _GEN_979;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_210 <= _GEN_6659;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_211 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_211 <= _GEN_980;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_211 <= _GEN_6660;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_212 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_212 <= _GEN_981;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_212 <= _GEN_6661;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_213 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_213 <= _GEN_982;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_213 <= _GEN_6662;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_214 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_214 <= _GEN_983;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_214 <= _GEN_6663;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_215 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_215 <= _GEN_984;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_215 <= _GEN_6664;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_216 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_216 <= _GEN_985;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_216 <= _GEN_6665;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_217 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_217 <= _GEN_986;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_217 <= _GEN_6666;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_218 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_218 <= _GEN_987;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_218 <= _GEN_6667;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_219 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_219 <= _GEN_988;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_219 <= _GEN_6668;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_220 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_220 <= _GEN_989;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_220 <= _GEN_6669;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_221 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_221 <= _GEN_990;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_221 <= _GEN_6670;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_222 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_222 <= _GEN_991;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_222 <= _GEN_6671;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_223 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_223 <= _GEN_992;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_223 <= _GEN_6672;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_224 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_224 <= _GEN_993;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_224 <= _GEN_6673;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_225 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_225 <= _GEN_994;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_225 <= _GEN_6674;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_226 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_226 <= _GEN_995;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_226 <= _GEN_6675;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_227 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_227 <= _GEN_996;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_227 <= _GEN_6676;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_228 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_228 <= _GEN_997;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_228 <= _GEN_6677;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_229 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_229 <= _GEN_998;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_229 <= _GEN_6678;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_230 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_230 <= _GEN_999;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_230 <= _GEN_6679;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_231 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_231 <= _GEN_1000;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_231 <= _GEN_6680;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_232 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_232 <= _GEN_1001;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_232 <= _GEN_6681;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_233 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_233 <= _GEN_1002;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_233 <= _GEN_6682;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_234 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_234 <= _GEN_1003;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_234 <= _GEN_6683;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_235 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_235 <= _GEN_1004;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_235 <= _GEN_6684;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_236 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_236 <= _GEN_1005;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_236 <= _GEN_6685;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_237 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_237 <= _GEN_1006;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_237 <= _GEN_6686;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_238 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_238 <= _GEN_1007;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_238 <= _GEN_6687;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_239 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_239 <= _GEN_1008;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_239 <= _GEN_6688;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_240 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_240 <= _GEN_1009;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_240 <= _GEN_6689;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_241 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_241 <= _GEN_1010;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_241 <= _GEN_6690;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_242 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_242 <= _GEN_1011;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_242 <= _GEN_6691;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_243 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_243 <= _GEN_1012;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_243 <= _GEN_6692;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_244 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_244 <= _GEN_1013;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_244 <= _GEN_6693;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_245 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_245 <= _GEN_1014;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_245 <= _GEN_6694;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_246 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_246 <= _GEN_1015;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_246 <= _GEN_6695;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_247 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_247 <= _GEN_1016;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_247 <= _GEN_6696;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_248 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_248 <= _GEN_1017;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_248 <= _GEN_6697;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_249 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_249 <= _GEN_1018;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_249 <= _GEN_6698;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_250 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_250 <= _GEN_1019;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_250 <= _GEN_6699;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_251 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_251 <= _GEN_1020;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_251 <= _GEN_6700;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_252 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_252 <= _GEN_1021;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_252 <= _GEN_6701;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_253 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_253 <= _GEN_1022;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_253 <= _GEN_6702;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_254 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_254 <= _GEN_1023;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_254 <= _GEN_6703;
      end
    end
    if (reset) begin // @[Dcache.scala 17:24]
      valid_255 <= 1'h0; // @[Dcache.scala 17:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          valid_255 <= _GEN_1024;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        valid_255 <= _GEN_6704;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_0 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_0 <= _GEN_1793;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_0 <= _GEN_6961;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_1 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_1 <= _GEN_1794;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_1 <= _GEN_6962;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_2 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_2 <= _GEN_1795;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_2 <= _GEN_6963;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_3 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_3 <= _GEN_1796;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_3 <= _GEN_6964;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_4 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_4 <= _GEN_1797;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_4 <= _GEN_6965;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_5 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_5 <= _GEN_1798;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_5 <= _GEN_6966;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_6 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_6 <= _GEN_1799;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_6 <= _GEN_6967;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_7 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_7 <= _GEN_1800;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_7 <= _GEN_6968;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_8 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_8 <= _GEN_1801;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_8 <= _GEN_6969;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_9 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_9 <= _GEN_1802;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_9 <= _GEN_6970;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_10 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_10 <= _GEN_1803;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_10 <= _GEN_6971;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_11 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_11 <= _GEN_1804;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_11 <= _GEN_6972;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_12 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_12 <= _GEN_1805;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_12 <= _GEN_6973;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_13 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_13 <= _GEN_1806;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_13 <= _GEN_6974;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_14 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_14 <= _GEN_1807;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_14 <= _GEN_6975;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_15 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_15 <= _GEN_1808;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_15 <= _GEN_6976;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_16 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_16 <= _GEN_1809;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_16 <= _GEN_6977;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_17 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_17 <= _GEN_1810;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_17 <= _GEN_6978;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_18 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_18 <= _GEN_1811;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_18 <= _GEN_6979;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_19 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_19 <= _GEN_1812;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_19 <= _GEN_6980;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_20 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_20 <= _GEN_1813;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_20 <= _GEN_6981;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_21 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_21 <= _GEN_1814;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_21 <= _GEN_6982;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_22 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_22 <= _GEN_1815;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_22 <= _GEN_6983;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_23 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_23 <= _GEN_1816;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_23 <= _GEN_6984;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_24 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_24 <= _GEN_1817;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_24 <= _GEN_6985;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_25 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_25 <= _GEN_1818;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_25 <= _GEN_6986;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_26 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_26 <= _GEN_1819;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_26 <= _GEN_6987;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_27 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_27 <= _GEN_1820;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_27 <= _GEN_6988;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_28 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_28 <= _GEN_1821;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_28 <= _GEN_6989;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_29 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_29 <= _GEN_1822;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_29 <= _GEN_6990;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_30 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_30 <= _GEN_1823;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_30 <= _GEN_6991;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_31 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_31 <= _GEN_1824;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_31 <= _GEN_6992;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_32 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_32 <= _GEN_1825;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_32 <= _GEN_6993;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_33 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_33 <= _GEN_1826;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_33 <= _GEN_6994;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_34 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_34 <= _GEN_1827;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_34 <= _GEN_6995;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_35 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_35 <= _GEN_1828;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_35 <= _GEN_6996;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_36 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_36 <= _GEN_1829;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_36 <= _GEN_6997;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_37 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_37 <= _GEN_1830;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_37 <= _GEN_6998;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_38 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_38 <= _GEN_1831;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_38 <= _GEN_6999;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_39 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_39 <= _GEN_1832;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_39 <= _GEN_7000;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_40 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_40 <= _GEN_1833;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_40 <= _GEN_7001;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_41 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_41 <= _GEN_1834;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_41 <= _GEN_7002;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_42 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_42 <= _GEN_1835;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_42 <= _GEN_7003;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_43 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_43 <= _GEN_1836;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_43 <= _GEN_7004;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_44 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_44 <= _GEN_1837;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_44 <= _GEN_7005;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_45 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_45 <= _GEN_1838;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_45 <= _GEN_7006;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_46 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_46 <= _GEN_1839;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_46 <= _GEN_7007;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_47 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_47 <= _GEN_1840;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_47 <= _GEN_7008;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_48 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_48 <= _GEN_1841;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_48 <= _GEN_7009;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_49 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_49 <= _GEN_1842;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_49 <= _GEN_7010;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_50 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_50 <= _GEN_1843;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_50 <= _GEN_7011;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_51 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_51 <= _GEN_1844;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_51 <= _GEN_7012;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_52 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_52 <= _GEN_1845;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_52 <= _GEN_7013;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_53 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_53 <= _GEN_1846;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_53 <= _GEN_7014;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_54 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_54 <= _GEN_1847;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_54 <= _GEN_7015;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_55 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_55 <= _GEN_1848;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_55 <= _GEN_7016;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_56 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_56 <= _GEN_1849;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_56 <= _GEN_7017;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_57 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_57 <= _GEN_1850;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_57 <= _GEN_7018;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_58 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_58 <= _GEN_1851;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_58 <= _GEN_7019;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_59 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_59 <= _GEN_1852;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_59 <= _GEN_7020;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_60 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_60 <= _GEN_1853;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_60 <= _GEN_7021;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_61 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_61 <= _GEN_1854;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_61 <= _GEN_7022;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_62 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_62 <= _GEN_1855;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_62 <= _GEN_7023;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_63 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_63 <= _GEN_1856;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_63 <= _GEN_7024;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_64 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_64 <= _GEN_1857;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_64 <= _GEN_7025;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_65 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_65 <= _GEN_1858;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_65 <= _GEN_7026;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_66 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_66 <= _GEN_1859;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_66 <= _GEN_7027;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_67 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_67 <= _GEN_1860;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_67 <= _GEN_7028;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_68 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_68 <= _GEN_1861;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_68 <= _GEN_7029;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_69 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_69 <= _GEN_1862;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_69 <= _GEN_7030;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_70 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_70 <= _GEN_1863;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_70 <= _GEN_7031;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_71 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_71 <= _GEN_1864;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_71 <= _GEN_7032;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_72 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_72 <= _GEN_1865;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_72 <= _GEN_7033;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_73 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_73 <= _GEN_1866;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_73 <= _GEN_7034;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_74 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_74 <= _GEN_1867;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_74 <= _GEN_7035;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_75 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_75 <= _GEN_1868;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_75 <= _GEN_7036;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_76 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_76 <= _GEN_1869;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_76 <= _GEN_7037;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_77 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_77 <= _GEN_1870;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_77 <= _GEN_7038;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_78 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_78 <= _GEN_1871;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_78 <= _GEN_7039;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_79 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_79 <= _GEN_1872;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_79 <= _GEN_7040;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_80 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_80 <= _GEN_1873;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_80 <= _GEN_7041;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_81 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_81 <= _GEN_1874;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_81 <= _GEN_7042;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_82 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_82 <= _GEN_1875;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_82 <= _GEN_7043;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_83 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_83 <= _GEN_1876;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_83 <= _GEN_7044;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_84 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_84 <= _GEN_1877;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_84 <= _GEN_7045;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_85 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_85 <= _GEN_1878;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_85 <= _GEN_7046;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_86 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_86 <= _GEN_1879;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_86 <= _GEN_7047;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_87 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_87 <= _GEN_1880;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_87 <= _GEN_7048;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_88 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_88 <= _GEN_1881;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_88 <= _GEN_7049;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_89 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_89 <= _GEN_1882;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_89 <= _GEN_7050;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_90 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_90 <= _GEN_1883;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_90 <= _GEN_7051;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_91 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_91 <= _GEN_1884;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_91 <= _GEN_7052;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_92 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_92 <= _GEN_1885;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_92 <= _GEN_7053;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_93 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_93 <= _GEN_1886;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_93 <= _GEN_7054;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_94 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_94 <= _GEN_1887;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_94 <= _GEN_7055;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_95 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_95 <= _GEN_1888;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_95 <= _GEN_7056;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_96 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_96 <= _GEN_1889;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_96 <= _GEN_7057;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_97 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_97 <= _GEN_1890;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_97 <= _GEN_7058;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_98 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_98 <= _GEN_1891;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_98 <= _GEN_7059;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_99 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_99 <= _GEN_1892;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_99 <= _GEN_7060;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_100 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_100 <= _GEN_1893;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_100 <= _GEN_7061;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_101 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_101 <= _GEN_1894;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_101 <= _GEN_7062;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_102 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_102 <= _GEN_1895;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_102 <= _GEN_7063;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_103 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_103 <= _GEN_1896;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_103 <= _GEN_7064;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_104 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_104 <= _GEN_1897;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_104 <= _GEN_7065;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_105 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_105 <= _GEN_1898;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_105 <= _GEN_7066;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_106 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_106 <= _GEN_1899;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_106 <= _GEN_7067;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_107 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_107 <= _GEN_1900;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_107 <= _GEN_7068;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_108 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_108 <= _GEN_1901;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_108 <= _GEN_7069;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_109 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_109 <= _GEN_1902;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_109 <= _GEN_7070;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_110 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_110 <= _GEN_1903;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_110 <= _GEN_7071;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_111 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_111 <= _GEN_1904;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_111 <= _GEN_7072;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_112 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_112 <= _GEN_1905;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_112 <= _GEN_7073;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_113 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_113 <= _GEN_1906;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_113 <= _GEN_7074;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_114 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_114 <= _GEN_1907;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_114 <= _GEN_7075;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_115 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_115 <= _GEN_1908;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_115 <= _GEN_7076;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_116 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_116 <= _GEN_1909;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_116 <= _GEN_7077;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_117 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_117 <= _GEN_1910;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_117 <= _GEN_7078;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_118 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_118 <= _GEN_1911;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_118 <= _GEN_7079;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_119 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_119 <= _GEN_1912;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_119 <= _GEN_7080;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_120 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_120 <= _GEN_1913;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_120 <= _GEN_7081;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_121 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_121 <= _GEN_1914;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_121 <= _GEN_7082;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_122 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_122 <= _GEN_1915;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_122 <= _GEN_7083;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_123 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_123 <= _GEN_1916;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_123 <= _GEN_7084;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_124 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_124 <= _GEN_1917;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_124 <= _GEN_7085;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_125 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_125 <= _GEN_1918;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_125 <= _GEN_7086;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_126 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_126 <= _GEN_1919;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_126 <= _GEN_7087;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_127 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_127 <= _GEN_1920;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_127 <= _GEN_7088;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_128 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_128 <= _GEN_1921;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_128 <= _GEN_7089;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_129 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_129 <= _GEN_1922;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_129 <= _GEN_7090;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_130 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_130 <= _GEN_1923;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_130 <= _GEN_7091;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_131 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_131 <= _GEN_1924;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_131 <= _GEN_7092;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_132 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_132 <= _GEN_1925;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_132 <= _GEN_7093;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_133 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_133 <= _GEN_1926;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_133 <= _GEN_7094;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_134 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_134 <= _GEN_1927;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_134 <= _GEN_7095;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_135 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_135 <= _GEN_1928;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_135 <= _GEN_7096;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_136 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_136 <= _GEN_1929;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_136 <= _GEN_7097;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_137 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_137 <= _GEN_1930;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_137 <= _GEN_7098;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_138 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_138 <= _GEN_1931;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_138 <= _GEN_7099;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_139 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_139 <= _GEN_1932;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_139 <= _GEN_7100;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_140 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_140 <= _GEN_1933;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_140 <= _GEN_7101;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_141 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_141 <= _GEN_1934;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_141 <= _GEN_7102;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_142 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_142 <= _GEN_1935;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_142 <= _GEN_7103;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_143 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_143 <= _GEN_1936;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_143 <= _GEN_7104;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_144 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_144 <= _GEN_1937;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_144 <= _GEN_7105;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_145 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_145 <= _GEN_1938;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_145 <= _GEN_7106;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_146 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_146 <= _GEN_1939;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_146 <= _GEN_7107;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_147 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_147 <= _GEN_1940;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_147 <= _GEN_7108;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_148 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_148 <= _GEN_1941;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_148 <= _GEN_7109;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_149 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_149 <= _GEN_1942;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_149 <= _GEN_7110;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_150 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_150 <= _GEN_1943;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_150 <= _GEN_7111;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_151 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_151 <= _GEN_1944;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_151 <= _GEN_7112;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_152 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_152 <= _GEN_1945;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_152 <= _GEN_7113;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_153 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_153 <= _GEN_1946;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_153 <= _GEN_7114;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_154 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_154 <= _GEN_1947;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_154 <= _GEN_7115;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_155 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_155 <= _GEN_1948;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_155 <= _GEN_7116;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_156 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_156 <= _GEN_1949;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_156 <= _GEN_7117;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_157 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_157 <= _GEN_1950;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_157 <= _GEN_7118;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_158 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_158 <= _GEN_1951;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_158 <= _GEN_7119;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_159 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_159 <= _GEN_1952;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_159 <= _GEN_7120;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_160 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_160 <= _GEN_1953;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_160 <= _GEN_7121;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_161 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_161 <= _GEN_1954;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_161 <= _GEN_7122;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_162 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_162 <= _GEN_1955;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_162 <= _GEN_7123;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_163 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_163 <= _GEN_1956;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_163 <= _GEN_7124;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_164 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_164 <= _GEN_1957;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_164 <= _GEN_7125;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_165 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_165 <= _GEN_1958;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_165 <= _GEN_7126;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_166 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_166 <= _GEN_1959;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_166 <= _GEN_7127;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_167 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_167 <= _GEN_1960;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_167 <= _GEN_7128;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_168 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_168 <= _GEN_1961;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_168 <= _GEN_7129;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_169 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_169 <= _GEN_1962;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_169 <= _GEN_7130;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_170 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_170 <= _GEN_1963;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_170 <= _GEN_7131;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_171 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_171 <= _GEN_1964;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_171 <= _GEN_7132;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_172 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_172 <= _GEN_1965;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_172 <= _GEN_7133;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_173 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_173 <= _GEN_1966;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_173 <= _GEN_7134;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_174 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_174 <= _GEN_1967;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_174 <= _GEN_7135;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_175 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_175 <= _GEN_1968;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_175 <= _GEN_7136;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_176 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_176 <= _GEN_1969;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_176 <= _GEN_7137;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_177 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_177 <= _GEN_1970;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_177 <= _GEN_7138;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_178 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_178 <= _GEN_1971;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_178 <= _GEN_7139;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_179 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_179 <= _GEN_1972;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_179 <= _GEN_7140;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_180 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_180 <= _GEN_1973;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_180 <= _GEN_7141;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_181 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_181 <= _GEN_1974;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_181 <= _GEN_7142;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_182 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_182 <= _GEN_1975;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_182 <= _GEN_7143;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_183 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_183 <= _GEN_1976;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_183 <= _GEN_7144;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_184 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_184 <= _GEN_1977;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_184 <= _GEN_7145;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_185 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_185 <= _GEN_1978;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_185 <= _GEN_7146;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_186 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_186 <= _GEN_1979;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_186 <= _GEN_7147;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_187 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_187 <= _GEN_1980;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_187 <= _GEN_7148;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_188 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_188 <= _GEN_1981;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_188 <= _GEN_7149;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_189 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_189 <= _GEN_1982;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_189 <= _GEN_7150;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_190 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_190 <= _GEN_1983;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_190 <= _GEN_7151;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_191 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_191 <= _GEN_1984;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_191 <= _GEN_7152;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_192 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_192 <= _GEN_1985;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_192 <= _GEN_7153;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_193 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_193 <= _GEN_1986;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_193 <= _GEN_7154;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_194 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_194 <= _GEN_1987;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_194 <= _GEN_7155;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_195 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_195 <= _GEN_1988;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_195 <= _GEN_7156;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_196 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_196 <= _GEN_1989;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_196 <= _GEN_7157;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_197 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_197 <= _GEN_1990;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_197 <= _GEN_7158;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_198 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_198 <= _GEN_1991;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_198 <= _GEN_7159;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_199 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_199 <= _GEN_1992;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_199 <= _GEN_7160;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_200 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_200 <= _GEN_1993;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_200 <= _GEN_7161;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_201 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_201 <= _GEN_1994;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_201 <= _GEN_7162;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_202 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_202 <= _GEN_1995;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_202 <= _GEN_7163;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_203 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_203 <= _GEN_1996;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_203 <= _GEN_7164;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_204 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_204 <= _GEN_1997;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_204 <= _GEN_7165;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_205 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_205 <= _GEN_1998;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_205 <= _GEN_7166;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_206 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_206 <= _GEN_1999;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_206 <= _GEN_7167;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_207 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_207 <= _GEN_2000;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_207 <= _GEN_7168;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_208 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_208 <= _GEN_2001;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_208 <= _GEN_7169;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_209 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_209 <= _GEN_2002;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_209 <= _GEN_7170;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_210 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_210 <= _GEN_2003;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_210 <= _GEN_7171;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_211 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_211 <= _GEN_2004;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_211 <= _GEN_7172;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_212 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_212 <= _GEN_2005;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_212 <= _GEN_7173;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_213 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_213 <= _GEN_2006;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_213 <= _GEN_7174;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_214 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_214 <= _GEN_2007;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_214 <= _GEN_7175;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_215 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_215 <= _GEN_2008;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_215 <= _GEN_7176;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_216 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_216 <= _GEN_2009;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_216 <= _GEN_7177;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_217 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_217 <= _GEN_2010;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_217 <= _GEN_7178;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_218 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_218 <= _GEN_2011;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_218 <= _GEN_7179;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_219 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_219 <= _GEN_2012;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_219 <= _GEN_7180;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_220 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_220 <= _GEN_2013;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_220 <= _GEN_7181;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_221 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_221 <= _GEN_2014;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_221 <= _GEN_7182;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_222 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_222 <= _GEN_2015;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_222 <= _GEN_7183;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_223 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_223 <= _GEN_2016;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_223 <= _GEN_7184;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_224 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_224 <= _GEN_2017;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_224 <= _GEN_7185;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_225 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_225 <= _GEN_2018;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_225 <= _GEN_7186;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_226 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_226 <= _GEN_2019;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_226 <= _GEN_7187;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_227 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_227 <= _GEN_2020;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_227 <= _GEN_7188;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_228 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_228 <= _GEN_2021;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_228 <= _GEN_7189;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_229 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_229 <= _GEN_2022;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_229 <= _GEN_7190;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_230 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_230 <= _GEN_2023;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_230 <= _GEN_7191;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_231 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_231 <= _GEN_2024;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_231 <= _GEN_7192;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_232 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_232 <= _GEN_2025;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_232 <= _GEN_7193;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_233 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_233 <= _GEN_2026;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_233 <= _GEN_7194;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_234 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_234 <= _GEN_2027;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_234 <= _GEN_7195;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_235 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_235 <= _GEN_2028;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_235 <= _GEN_7196;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_236 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_236 <= _GEN_2029;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_236 <= _GEN_7197;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_237 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_237 <= _GEN_2030;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_237 <= _GEN_7198;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_238 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_238 <= _GEN_2031;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_238 <= _GEN_7199;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_239 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_239 <= _GEN_2032;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_239 <= _GEN_7200;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_240 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_240 <= _GEN_2033;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_240 <= _GEN_7201;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_241 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_241 <= _GEN_2034;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_241 <= _GEN_7202;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_242 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_242 <= _GEN_2035;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_242 <= _GEN_7203;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_243 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_243 <= _GEN_2036;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_243 <= _GEN_7204;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_244 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_244 <= _GEN_2037;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_244 <= _GEN_7205;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_245 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_245 <= _GEN_2038;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_245 <= _GEN_7206;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_246 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_246 <= _GEN_2039;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_246 <= _GEN_7207;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_247 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_247 <= _GEN_2040;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_247 <= _GEN_7208;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_248 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_248 <= _GEN_2041;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_248 <= _GEN_7209;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_249 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_249 <= _GEN_2042;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_249 <= _GEN_7210;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_250 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_250 <= _GEN_2043;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_250 <= _GEN_7211;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_251 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_251 <= _GEN_2044;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_251 <= _GEN_7212;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_252 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_252 <= _GEN_2045;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_252 <= _GEN_7213;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_253 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_253 <= _GEN_2046;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_253 <= _GEN_7214;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_254 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_254 <= _GEN_2047;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_254 <= _GEN_7215;
      end
    end
    if (reset) begin // @[Dcache.scala 18:24]
      dirty_255 <= 1'h0; // @[Dcache.scala 18:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          dirty_255 <= _GEN_2048;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        dirty_255 <= _GEN_7216;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_0 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_0 <= _GEN_1281;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_0 <= _GEN_7217;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_1 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_1 <= _GEN_1282;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_1 <= _GEN_7218;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_2 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_2 <= _GEN_1283;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_2 <= _GEN_7219;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_3 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_3 <= _GEN_1284;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_3 <= _GEN_7220;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_4 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_4 <= _GEN_1285;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_4 <= _GEN_7221;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_5 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_5 <= _GEN_1286;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_5 <= _GEN_7222;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_6 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_6 <= _GEN_1287;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_6 <= _GEN_7223;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_7 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_7 <= _GEN_1288;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_7 <= _GEN_7224;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_8 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_8 <= _GEN_1289;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_8 <= _GEN_7225;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_9 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_9 <= _GEN_1290;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_9 <= _GEN_7226;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_10 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_10 <= _GEN_1291;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_10 <= _GEN_7227;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_11 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_11 <= _GEN_1292;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_11 <= _GEN_7228;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_12 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_12 <= _GEN_1293;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_12 <= _GEN_7229;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_13 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_13 <= _GEN_1294;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_13 <= _GEN_7230;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_14 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_14 <= _GEN_1295;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_14 <= _GEN_7231;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_15 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_15 <= _GEN_1296;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_15 <= _GEN_7232;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_16 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_16 <= _GEN_1297;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_16 <= _GEN_7233;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_17 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_17 <= _GEN_1298;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_17 <= _GEN_7234;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_18 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_18 <= _GEN_1299;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_18 <= _GEN_7235;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_19 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_19 <= _GEN_1300;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_19 <= _GEN_7236;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_20 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_20 <= _GEN_1301;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_20 <= _GEN_7237;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_21 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_21 <= _GEN_1302;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_21 <= _GEN_7238;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_22 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_22 <= _GEN_1303;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_22 <= _GEN_7239;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_23 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_23 <= _GEN_1304;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_23 <= _GEN_7240;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_24 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_24 <= _GEN_1305;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_24 <= _GEN_7241;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_25 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_25 <= _GEN_1306;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_25 <= _GEN_7242;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_26 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_26 <= _GEN_1307;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_26 <= _GEN_7243;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_27 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_27 <= _GEN_1308;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_27 <= _GEN_7244;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_28 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_28 <= _GEN_1309;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_28 <= _GEN_7245;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_29 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_29 <= _GEN_1310;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_29 <= _GEN_7246;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_30 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_30 <= _GEN_1311;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_30 <= _GEN_7247;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_31 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_31 <= _GEN_1312;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_31 <= _GEN_7248;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_32 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_32 <= _GEN_1313;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_32 <= _GEN_7249;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_33 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_33 <= _GEN_1314;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_33 <= _GEN_7250;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_34 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_34 <= _GEN_1315;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_34 <= _GEN_7251;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_35 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_35 <= _GEN_1316;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_35 <= _GEN_7252;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_36 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_36 <= _GEN_1317;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_36 <= _GEN_7253;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_37 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_37 <= _GEN_1318;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_37 <= _GEN_7254;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_38 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_38 <= _GEN_1319;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_38 <= _GEN_7255;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_39 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_39 <= _GEN_1320;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_39 <= _GEN_7256;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_40 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_40 <= _GEN_1321;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_40 <= _GEN_7257;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_41 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_41 <= _GEN_1322;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_41 <= _GEN_7258;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_42 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_42 <= _GEN_1323;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_42 <= _GEN_7259;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_43 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_43 <= _GEN_1324;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_43 <= _GEN_7260;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_44 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_44 <= _GEN_1325;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_44 <= _GEN_7261;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_45 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_45 <= _GEN_1326;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_45 <= _GEN_7262;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_46 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_46 <= _GEN_1327;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_46 <= _GEN_7263;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_47 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_47 <= _GEN_1328;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_47 <= _GEN_7264;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_48 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_48 <= _GEN_1329;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_48 <= _GEN_7265;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_49 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_49 <= _GEN_1330;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_49 <= _GEN_7266;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_50 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_50 <= _GEN_1331;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_50 <= _GEN_7267;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_51 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_51 <= _GEN_1332;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_51 <= _GEN_7268;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_52 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_52 <= _GEN_1333;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_52 <= _GEN_7269;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_53 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_53 <= _GEN_1334;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_53 <= _GEN_7270;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_54 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_54 <= _GEN_1335;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_54 <= _GEN_7271;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_55 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_55 <= _GEN_1336;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_55 <= _GEN_7272;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_56 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_56 <= _GEN_1337;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_56 <= _GEN_7273;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_57 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_57 <= _GEN_1338;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_57 <= _GEN_7274;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_58 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_58 <= _GEN_1339;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_58 <= _GEN_7275;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_59 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_59 <= _GEN_1340;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_59 <= _GEN_7276;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_60 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_60 <= _GEN_1341;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_60 <= _GEN_7277;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_61 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_61 <= _GEN_1342;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_61 <= _GEN_7278;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_62 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_62 <= _GEN_1343;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_62 <= _GEN_7279;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_63 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_63 <= _GEN_1344;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_63 <= _GEN_7280;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_64 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_64 <= _GEN_1345;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_64 <= _GEN_7281;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_65 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_65 <= _GEN_1346;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_65 <= _GEN_7282;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_66 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_66 <= _GEN_1347;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_66 <= _GEN_7283;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_67 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_67 <= _GEN_1348;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_67 <= _GEN_7284;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_68 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_68 <= _GEN_1349;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_68 <= _GEN_7285;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_69 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_69 <= _GEN_1350;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_69 <= _GEN_7286;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_70 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_70 <= _GEN_1351;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_70 <= _GEN_7287;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_71 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_71 <= _GEN_1352;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_71 <= _GEN_7288;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_72 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_72 <= _GEN_1353;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_72 <= _GEN_7289;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_73 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_73 <= _GEN_1354;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_73 <= _GEN_7290;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_74 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_74 <= _GEN_1355;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_74 <= _GEN_7291;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_75 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_75 <= _GEN_1356;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_75 <= _GEN_7292;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_76 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_76 <= _GEN_1357;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_76 <= _GEN_7293;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_77 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_77 <= _GEN_1358;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_77 <= _GEN_7294;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_78 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_78 <= _GEN_1359;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_78 <= _GEN_7295;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_79 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_79 <= _GEN_1360;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_79 <= _GEN_7296;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_80 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_80 <= _GEN_1361;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_80 <= _GEN_7297;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_81 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_81 <= _GEN_1362;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_81 <= _GEN_7298;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_82 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_82 <= _GEN_1363;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_82 <= _GEN_7299;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_83 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_83 <= _GEN_1364;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_83 <= _GEN_7300;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_84 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_84 <= _GEN_1365;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_84 <= _GEN_7301;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_85 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_85 <= _GEN_1366;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_85 <= _GEN_7302;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_86 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_86 <= _GEN_1367;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_86 <= _GEN_7303;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_87 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_87 <= _GEN_1368;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_87 <= _GEN_7304;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_88 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_88 <= _GEN_1369;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_88 <= _GEN_7305;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_89 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_89 <= _GEN_1370;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_89 <= _GEN_7306;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_90 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_90 <= _GEN_1371;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_90 <= _GEN_7307;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_91 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_91 <= _GEN_1372;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_91 <= _GEN_7308;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_92 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_92 <= _GEN_1373;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_92 <= _GEN_7309;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_93 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_93 <= _GEN_1374;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_93 <= _GEN_7310;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_94 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_94 <= _GEN_1375;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_94 <= _GEN_7311;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_95 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_95 <= _GEN_1376;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_95 <= _GEN_7312;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_96 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_96 <= _GEN_1377;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_96 <= _GEN_7313;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_97 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_97 <= _GEN_1378;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_97 <= _GEN_7314;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_98 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_98 <= _GEN_1379;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_98 <= _GEN_7315;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_99 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_99 <= _GEN_1380;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_99 <= _GEN_7316;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_100 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_100 <= _GEN_1381;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_100 <= _GEN_7317;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_101 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_101 <= _GEN_1382;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_101 <= _GEN_7318;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_102 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_102 <= _GEN_1383;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_102 <= _GEN_7319;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_103 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_103 <= _GEN_1384;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_103 <= _GEN_7320;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_104 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_104 <= _GEN_1385;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_104 <= _GEN_7321;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_105 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_105 <= _GEN_1386;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_105 <= _GEN_7322;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_106 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_106 <= _GEN_1387;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_106 <= _GEN_7323;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_107 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_107 <= _GEN_1388;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_107 <= _GEN_7324;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_108 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_108 <= _GEN_1389;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_108 <= _GEN_7325;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_109 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_109 <= _GEN_1390;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_109 <= _GEN_7326;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_110 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_110 <= _GEN_1391;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_110 <= _GEN_7327;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_111 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_111 <= _GEN_1392;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_111 <= _GEN_7328;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_112 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_112 <= _GEN_1393;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_112 <= _GEN_7329;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_113 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_113 <= _GEN_1394;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_113 <= _GEN_7330;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_114 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_114 <= _GEN_1395;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_114 <= _GEN_7331;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_115 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_115 <= _GEN_1396;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_115 <= _GEN_7332;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_116 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_116 <= _GEN_1397;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_116 <= _GEN_7333;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_117 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_117 <= _GEN_1398;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_117 <= _GEN_7334;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_118 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_118 <= _GEN_1399;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_118 <= _GEN_7335;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_119 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_119 <= _GEN_1400;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_119 <= _GEN_7336;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_120 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_120 <= _GEN_1401;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_120 <= _GEN_7337;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_121 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_121 <= _GEN_1402;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_121 <= _GEN_7338;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_122 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_122 <= _GEN_1403;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_122 <= _GEN_7339;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_123 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_123 <= _GEN_1404;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_123 <= _GEN_7340;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_124 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_124 <= _GEN_1405;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_124 <= _GEN_7341;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_125 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_125 <= _GEN_1406;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_125 <= _GEN_7342;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_126 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_126 <= _GEN_1407;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_126 <= _GEN_7343;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_127 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_127 <= _GEN_1408;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_127 <= _GEN_7344;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_128 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_128 <= _GEN_1409;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_128 <= _GEN_7345;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_129 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_129 <= _GEN_1410;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_129 <= _GEN_7346;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_130 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_130 <= _GEN_1411;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_130 <= _GEN_7347;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_131 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_131 <= _GEN_1412;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_131 <= _GEN_7348;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_132 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_132 <= _GEN_1413;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_132 <= _GEN_7349;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_133 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_133 <= _GEN_1414;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_133 <= _GEN_7350;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_134 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_134 <= _GEN_1415;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_134 <= _GEN_7351;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_135 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_135 <= _GEN_1416;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_135 <= _GEN_7352;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_136 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_136 <= _GEN_1417;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_136 <= _GEN_7353;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_137 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_137 <= _GEN_1418;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_137 <= _GEN_7354;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_138 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_138 <= _GEN_1419;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_138 <= _GEN_7355;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_139 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_139 <= _GEN_1420;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_139 <= _GEN_7356;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_140 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_140 <= _GEN_1421;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_140 <= _GEN_7357;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_141 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_141 <= _GEN_1422;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_141 <= _GEN_7358;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_142 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_142 <= _GEN_1423;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_142 <= _GEN_7359;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_143 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_143 <= _GEN_1424;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_143 <= _GEN_7360;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_144 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_144 <= _GEN_1425;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_144 <= _GEN_7361;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_145 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_145 <= _GEN_1426;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_145 <= _GEN_7362;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_146 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_146 <= _GEN_1427;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_146 <= _GEN_7363;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_147 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_147 <= _GEN_1428;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_147 <= _GEN_7364;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_148 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_148 <= _GEN_1429;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_148 <= _GEN_7365;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_149 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_149 <= _GEN_1430;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_149 <= _GEN_7366;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_150 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_150 <= _GEN_1431;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_150 <= _GEN_7367;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_151 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_151 <= _GEN_1432;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_151 <= _GEN_7368;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_152 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_152 <= _GEN_1433;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_152 <= _GEN_7369;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_153 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_153 <= _GEN_1434;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_153 <= _GEN_7370;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_154 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_154 <= _GEN_1435;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_154 <= _GEN_7371;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_155 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_155 <= _GEN_1436;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_155 <= _GEN_7372;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_156 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_156 <= _GEN_1437;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_156 <= _GEN_7373;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_157 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_157 <= _GEN_1438;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_157 <= _GEN_7374;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_158 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_158 <= _GEN_1439;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_158 <= _GEN_7375;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_159 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_159 <= _GEN_1440;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_159 <= _GEN_7376;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_160 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_160 <= _GEN_1441;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_160 <= _GEN_7377;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_161 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_161 <= _GEN_1442;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_161 <= _GEN_7378;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_162 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_162 <= _GEN_1443;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_162 <= _GEN_7379;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_163 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_163 <= _GEN_1444;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_163 <= _GEN_7380;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_164 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_164 <= _GEN_1445;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_164 <= _GEN_7381;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_165 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_165 <= _GEN_1446;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_165 <= _GEN_7382;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_166 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_166 <= _GEN_1447;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_166 <= _GEN_7383;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_167 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_167 <= _GEN_1448;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_167 <= _GEN_7384;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_168 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_168 <= _GEN_1449;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_168 <= _GEN_7385;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_169 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_169 <= _GEN_1450;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_169 <= _GEN_7386;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_170 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_170 <= _GEN_1451;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_170 <= _GEN_7387;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_171 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_171 <= _GEN_1452;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_171 <= _GEN_7388;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_172 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_172 <= _GEN_1453;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_172 <= _GEN_7389;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_173 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_173 <= _GEN_1454;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_173 <= _GEN_7390;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_174 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_174 <= _GEN_1455;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_174 <= _GEN_7391;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_175 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_175 <= _GEN_1456;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_175 <= _GEN_7392;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_176 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_176 <= _GEN_1457;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_176 <= _GEN_7393;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_177 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_177 <= _GEN_1458;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_177 <= _GEN_7394;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_178 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_178 <= _GEN_1459;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_178 <= _GEN_7395;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_179 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_179 <= _GEN_1460;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_179 <= _GEN_7396;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_180 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_180 <= _GEN_1461;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_180 <= _GEN_7397;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_181 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_181 <= _GEN_1462;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_181 <= _GEN_7398;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_182 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_182 <= _GEN_1463;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_182 <= _GEN_7399;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_183 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_183 <= _GEN_1464;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_183 <= _GEN_7400;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_184 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_184 <= _GEN_1465;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_184 <= _GEN_7401;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_185 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_185 <= _GEN_1466;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_185 <= _GEN_7402;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_186 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_186 <= _GEN_1467;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_186 <= _GEN_7403;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_187 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_187 <= _GEN_1468;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_187 <= _GEN_7404;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_188 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_188 <= _GEN_1469;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_188 <= _GEN_7405;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_189 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_189 <= _GEN_1470;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_189 <= _GEN_7406;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_190 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_190 <= _GEN_1471;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_190 <= _GEN_7407;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_191 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_191 <= _GEN_1472;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_191 <= _GEN_7408;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_192 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_192 <= _GEN_1473;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_192 <= _GEN_7409;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_193 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_193 <= _GEN_1474;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_193 <= _GEN_7410;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_194 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_194 <= _GEN_1475;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_194 <= _GEN_7411;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_195 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_195 <= _GEN_1476;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_195 <= _GEN_7412;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_196 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_196 <= _GEN_1477;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_196 <= _GEN_7413;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_197 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_197 <= _GEN_1478;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_197 <= _GEN_7414;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_198 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_198 <= _GEN_1479;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_198 <= _GEN_7415;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_199 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_199 <= _GEN_1480;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_199 <= _GEN_7416;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_200 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_200 <= _GEN_1481;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_200 <= _GEN_7417;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_201 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_201 <= _GEN_1482;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_201 <= _GEN_7418;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_202 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_202 <= _GEN_1483;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_202 <= _GEN_7419;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_203 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_203 <= _GEN_1484;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_203 <= _GEN_7420;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_204 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_204 <= _GEN_1485;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_204 <= _GEN_7421;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_205 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_205 <= _GEN_1486;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_205 <= _GEN_7422;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_206 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_206 <= _GEN_1487;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_206 <= _GEN_7423;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_207 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_207 <= _GEN_1488;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_207 <= _GEN_7424;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_208 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_208 <= _GEN_1489;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_208 <= _GEN_7425;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_209 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_209 <= _GEN_1490;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_209 <= _GEN_7426;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_210 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_210 <= _GEN_1491;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_210 <= _GEN_7427;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_211 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_211 <= _GEN_1492;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_211 <= _GEN_7428;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_212 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_212 <= _GEN_1493;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_212 <= _GEN_7429;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_213 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_213 <= _GEN_1494;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_213 <= _GEN_7430;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_214 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_214 <= _GEN_1495;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_214 <= _GEN_7431;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_215 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_215 <= _GEN_1496;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_215 <= _GEN_7432;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_216 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_216 <= _GEN_1497;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_216 <= _GEN_7433;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_217 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_217 <= _GEN_1498;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_217 <= _GEN_7434;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_218 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_218 <= _GEN_1499;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_218 <= _GEN_7435;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_219 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_219 <= _GEN_1500;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_219 <= _GEN_7436;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_220 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_220 <= _GEN_1501;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_220 <= _GEN_7437;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_221 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_221 <= _GEN_1502;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_221 <= _GEN_7438;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_222 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_222 <= _GEN_1503;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_222 <= _GEN_7439;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_223 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_223 <= _GEN_1504;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_223 <= _GEN_7440;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_224 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_224 <= _GEN_1505;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_224 <= _GEN_7441;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_225 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_225 <= _GEN_1506;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_225 <= _GEN_7442;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_226 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_226 <= _GEN_1507;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_226 <= _GEN_7443;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_227 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_227 <= _GEN_1508;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_227 <= _GEN_7444;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_228 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_228 <= _GEN_1509;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_228 <= _GEN_7445;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_229 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_229 <= _GEN_1510;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_229 <= _GEN_7446;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_230 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_230 <= _GEN_1511;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_230 <= _GEN_7447;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_231 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_231 <= _GEN_1512;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_231 <= _GEN_7448;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_232 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_232 <= _GEN_1513;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_232 <= _GEN_7449;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_233 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_233 <= _GEN_1514;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_233 <= _GEN_7450;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_234 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_234 <= _GEN_1515;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_234 <= _GEN_7451;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_235 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_235 <= _GEN_1516;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_235 <= _GEN_7452;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_236 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_236 <= _GEN_1517;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_236 <= _GEN_7453;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_237 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_237 <= _GEN_1518;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_237 <= _GEN_7454;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_238 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_238 <= _GEN_1519;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_238 <= _GEN_7455;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_239 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_239 <= _GEN_1520;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_239 <= _GEN_7456;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_240 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_240 <= _GEN_1521;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_240 <= _GEN_7457;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_241 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_241 <= _GEN_1522;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_241 <= _GEN_7458;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_242 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_242 <= _GEN_1523;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_242 <= _GEN_7459;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_243 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_243 <= _GEN_1524;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_243 <= _GEN_7460;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_244 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_244 <= _GEN_1525;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_244 <= _GEN_7461;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_245 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_245 <= _GEN_1526;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_245 <= _GEN_7462;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_246 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_246 <= _GEN_1527;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_246 <= _GEN_7463;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_247 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_247 <= _GEN_1528;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_247 <= _GEN_7464;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_248 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_248 <= _GEN_1529;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_248 <= _GEN_7465;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_249 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_249 <= _GEN_1530;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_249 <= _GEN_7466;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_250 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_250 <= _GEN_1531;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_250 <= _GEN_7467;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_251 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_251 <= _GEN_1532;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_251 <= _GEN_7468;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_252 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_252 <= _GEN_1533;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_252 <= _GEN_7469;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_253 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_253 <= _GEN_1534;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_253 <= _GEN_7470;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_254 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_254 <= _GEN_1535;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_254 <= _GEN_7471;
      end
    end
    if (reset) begin // @[Dcache.scala 19:24]
      offset_255 <= 4'h0; // @[Dcache.scala 19:24]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          offset_255 <= _GEN_1536;
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        offset_255 <= _GEN_7472;
      end
    end
    if (reset) begin // @[Dcache.scala 26:22]
      state <= 3'h0; // @[Dcache.scala 26:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_dmem_data_valid) begin // @[Dcache.scala 125:28]
        state <= 3'h1; // @[Dcache.scala 126:15]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (cache_hit) begin // @[Dcache.scala 131:24]
        state <= 3'h0; // @[Dcache.scala 142:27]
      end else begin
        state <= _GEN_2049;
      end
    end else if (_T_3) begin // @[Conditional.scala 39:67]
      state <= _GEN_3335;
    end else begin
      state <= _GEN_6437;
    end
    if (reset) begin // @[Dcache.scala 46:28]
      data_ready <= 1'h0; // @[Dcache.scala 46:28]
    end else if (_T) begin // @[Conditional.scala 40:58]
      data_ready <= 1'h0; // @[Dcache.scala 123:18]
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      data_ready <= _GEN_2818;
    end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
      data_ready <= _GEN_6448;
    end
    if (reset) begin // @[Dcache.scala 116:28]
      cache_fill <= 1'h0; // @[Dcache.scala 116:28]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_1)) begin // @[Conditional.scala 39:67]
        if (!(_T_3)) begin // @[Conditional.scala 39:67]
          cache_fill <= _GEN_6444;
        end
      end
    end
    if (reset) begin // @[Dcache.scala 117:28]
      cache_wen <= 1'h0; // @[Dcache.scala 117:28]
    end else if (_T) begin // @[Conditional.scala 40:58]
      cache_wen <= 1'h0; // @[Dcache.scala 124:18]
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (cache_hit) begin // @[Dcache.scala 131:24]
        cache_wen <= io_dmem_data_req; // @[Dcache.scala 136:27]
      end
    end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
      cache_wen <= _GEN_6445;
    end
    if (reset) begin // @[Dcache.scala 118:28]
      cache_wdata <= 128'h0; // @[Dcache.scala 118:28]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          cache_wdata <= _cache_wdata_T_3; // @[Dcache.scala 137:27]
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        cache_wdata <= _GEN_6446;
      end
    end
    if (reset) begin // @[Dcache.scala 119:28]
      cache_strb <= 128'h0; // @[Dcache.scala 119:28]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (cache_hit) begin // @[Dcache.scala 131:24]
          cache_strb <= _cache_strb_T_3; // @[Dcache.scala 138:27]
        end
      end else if (!(_T_3)) begin // @[Conditional.scala 39:67]
        cache_strb <= _GEN_6447;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_0 = _RAND_0[19:0];
  _RAND_1 = {1{`RANDOM}};
  tag_1 = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  tag_2 = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  tag_3 = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  tag_4 = _RAND_4[19:0];
  _RAND_5 = {1{`RANDOM}};
  tag_5 = _RAND_5[19:0];
  _RAND_6 = {1{`RANDOM}};
  tag_6 = _RAND_6[19:0];
  _RAND_7 = {1{`RANDOM}};
  tag_7 = _RAND_7[19:0];
  _RAND_8 = {1{`RANDOM}};
  tag_8 = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  tag_9 = _RAND_9[19:0];
  _RAND_10 = {1{`RANDOM}};
  tag_10 = _RAND_10[19:0];
  _RAND_11 = {1{`RANDOM}};
  tag_11 = _RAND_11[19:0];
  _RAND_12 = {1{`RANDOM}};
  tag_12 = _RAND_12[19:0];
  _RAND_13 = {1{`RANDOM}};
  tag_13 = _RAND_13[19:0];
  _RAND_14 = {1{`RANDOM}};
  tag_14 = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  tag_15 = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  tag_16 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  tag_17 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  tag_18 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  tag_19 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  tag_20 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  tag_21 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  tag_22 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  tag_23 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  tag_24 = _RAND_24[19:0];
  _RAND_25 = {1{`RANDOM}};
  tag_25 = _RAND_25[19:0];
  _RAND_26 = {1{`RANDOM}};
  tag_26 = _RAND_26[19:0];
  _RAND_27 = {1{`RANDOM}};
  tag_27 = _RAND_27[19:0];
  _RAND_28 = {1{`RANDOM}};
  tag_28 = _RAND_28[19:0];
  _RAND_29 = {1{`RANDOM}};
  tag_29 = _RAND_29[19:0];
  _RAND_30 = {1{`RANDOM}};
  tag_30 = _RAND_30[19:0];
  _RAND_31 = {1{`RANDOM}};
  tag_31 = _RAND_31[19:0];
  _RAND_32 = {1{`RANDOM}};
  tag_32 = _RAND_32[19:0];
  _RAND_33 = {1{`RANDOM}};
  tag_33 = _RAND_33[19:0];
  _RAND_34 = {1{`RANDOM}};
  tag_34 = _RAND_34[19:0];
  _RAND_35 = {1{`RANDOM}};
  tag_35 = _RAND_35[19:0];
  _RAND_36 = {1{`RANDOM}};
  tag_36 = _RAND_36[19:0];
  _RAND_37 = {1{`RANDOM}};
  tag_37 = _RAND_37[19:0];
  _RAND_38 = {1{`RANDOM}};
  tag_38 = _RAND_38[19:0];
  _RAND_39 = {1{`RANDOM}};
  tag_39 = _RAND_39[19:0];
  _RAND_40 = {1{`RANDOM}};
  tag_40 = _RAND_40[19:0];
  _RAND_41 = {1{`RANDOM}};
  tag_41 = _RAND_41[19:0];
  _RAND_42 = {1{`RANDOM}};
  tag_42 = _RAND_42[19:0];
  _RAND_43 = {1{`RANDOM}};
  tag_43 = _RAND_43[19:0];
  _RAND_44 = {1{`RANDOM}};
  tag_44 = _RAND_44[19:0];
  _RAND_45 = {1{`RANDOM}};
  tag_45 = _RAND_45[19:0];
  _RAND_46 = {1{`RANDOM}};
  tag_46 = _RAND_46[19:0];
  _RAND_47 = {1{`RANDOM}};
  tag_47 = _RAND_47[19:0];
  _RAND_48 = {1{`RANDOM}};
  tag_48 = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  tag_49 = _RAND_49[19:0];
  _RAND_50 = {1{`RANDOM}};
  tag_50 = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  tag_51 = _RAND_51[19:0];
  _RAND_52 = {1{`RANDOM}};
  tag_52 = _RAND_52[19:0];
  _RAND_53 = {1{`RANDOM}};
  tag_53 = _RAND_53[19:0];
  _RAND_54 = {1{`RANDOM}};
  tag_54 = _RAND_54[19:0];
  _RAND_55 = {1{`RANDOM}};
  tag_55 = _RAND_55[19:0];
  _RAND_56 = {1{`RANDOM}};
  tag_56 = _RAND_56[19:0];
  _RAND_57 = {1{`RANDOM}};
  tag_57 = _RAND_57[19:0];
  _RAND_58 = {1{`RANDOM}};
  tag_58 = _RAND_58[19:0];
  _RAND_59 = {1{`RANDOM}};
  tag_59 = _RAND_59[19:0];
  _RAND_60 = {1{`RANDOM}};
  tag_60 = _RAND_60[19:0];
  _RAND_61 = {1{`RANDOM}};
  tag_61 = _RAND_61[19:0];
  _RAND_62 = {1{`RANDOM}};
  tag_62 = _RAND_62[19:0];
  _RAND_63 = {1{`RANDOM}};
  tag_63 = _RAND_63[19:0];
  _RAND_64 = {1{`RANDOM}};
  tag_64 = _RAND_64[19:0];
  _RAND_65 = {1{`RANDOM}};
  tag_65 = _RAND_65[19:0];
  _RAND_66 = {1{`RANDOM}};
  tag_66 = _RAND_66[19:0];
  _RAND_67 = {1{`RANDOM}};
  tag_67 = _RAND_67[19:0];
  _RAND_68 = {1{`RANDOM}};
  tag_68 = _RAND_68[19:0];
  _RAND_69 = {1{`RANDOM}};
  tag_69 = _RAND_69[19:0];
  _RAND_70 = {1{`RANDOM}};
  tag_70 = _RAND_70[19:0];
  _RAND_71 = {1{`RANDOM}};
  tag_71 = _RAND_71[19:0];
  _RAND_72 = {1{`RANDOM}};
  tag_72 = _RAND_72[19:0];
  _RAND_73 = {1{`RANDOM}};
  tag_73 = _RAND_73[19:0];
  _RAND_74 = {1{`RANDOM}};
  tag_74 = _RAND_74[19:0];
  _RAND_75 = {1{`RANDOM}};
  tag_75 = _RAND_75[19:0];
  _RAND_76 = {1{`RANDOM}};
  tag_76 = _RAND_76[19:0];
  _RAND_77 = {1{`RANDOM}};
  tag_77 = _RAND_77[19:0];
  _RAND_78 = {1{`RANDOM}};
  tag_78 = _RAND_78[19:0];
  _RAND_79 = {1{`RANDOM}};
  tag_79 = _RAND_79[19:0];
  _RAND_80 = {1{`RANDOM}};
  tag_80 = _RAND_80[19:0];
  _RAND_81 = {1{`RANDOM}};
  tag_81 = _RAND_81[19:0];
  _RAND_82 = {1{`RANDOM}};
  tag_82 = _RAND_82[19:0];
  _RAND_83 = {1{`RANDOM}};
  tag_83 = _RAND_83[19:0];
  _RAND_84 = {1{`RANDOM}};
  tag_84 = _RAND_84[19:0];
  _RAND_85 = {1{`RANDOM}};
  tag_85 = _RAND_85[19:0];
  _RAND_86 = {1{`RANDOM}};
  tag_86 = _RAND_86[19:0];
  _RAND_87 = {1{`RANDOM}};
  tag_87 = _RAND_87[19:0];
  _RAND_88 = {1{`RANDOM}};
  tag_88 = _RAND_88[19:0];
  _RAND_89 = {1{`RANDOM}};
  tag_89 = _RAND_89[19:0];
  _RAND_90 = {1{`RANDOM}};
  tag_90 = _RAND_90[19:0];
  _RAND_91 = {1{`RANDOM}};
  tag_91 = _RAND_91[19:0];
  _RAND_92 = {1{`RANDOM}};
  tag_92 = _RAND_92[19:0];
  _RAND_93 = {1{`RANDOM}};
  tag_93 = _RAND_93[19:0];
  _RAND_94 = {1{`RANDOM}};
  tag_94 = _RAND_94[19:0];
  _RAND_95 = {1{`RANDOM}};
  tag_95 = _RAND_95[19:0];
  _RAND_96 = {1{`RANDOM}};
  tag_96 = _RAND_96[19:0];
  _RAND_97 = {1{`RANDOM}};
  tag_97 = _RAND_97[19:0];
  _RAND_98 = {1{`RANDOM}};
  tag_98 = _RAND_98[19:0];
  _RAND_99 = {1{`RANDOM}};
  tag_99 = _RAND_99[19:0];
  _RAND_100 = {1{`RANDOM}};
  tag_100 = _RAND_100[19:0];
  _RAND_101 = {1{`RANDOM}};
  tag_101 = _RAND_101[19:0];
  _RAND_102 = {1{`RANDOM}};
  tag_102 = _RAND_102[19:0];
  _RAND_103 = {1{`RANDOM}};
  tag_103 = _RAND_103[19:0];
  _RAND_104 = {1{`RANDOM}};
  tag_104 = _RAND_104[19:0];
  _RAND_105 = {1{`RANDOM}};
  tag_105 = _RAND_105[19:0];
  _RAND_106 = {1{`RANDOM}};
  tag_106 = _RAND_106[19:0];
  _RAND_107 = {1{`RANDOM}};
  tag_107 = _RAND_107[19:0];
  _RAND_108 = {1{`RANDOM}};
  tag_108 = _RAND_108[19:0];
  _RAND_109 = {1{`RANDOM}};
  tag_109 = _RAND_109[19:0];
  _RAND_110 = {1{`RANDOM}};
  tag_110 = _RAND_110[19:0];
  _RAND_111 = {1{`RANDOM}};
  tag_111 = _RAND_111[19:0];
  _RAND_112 = {1{`RANDOM}};
  tag_112 = _RAND_112[19:0];
  _RAND_113 = {1{`RANDOM}};
  tag_113 = _RAND_113[19:0];
  _RAND_114 = {1{`RANDOM}};
  tag_114 = _RAND_114[19:0];
  _RAND_115 = {1{`RANDOM}};
  tag_115 = _RAND_115[19:0];
  _RAND_116 = {1{`RANDOM}};
  tag_116 = _RAND_116[19:0];
  _RAND_117 = {1{`RANDOM}};
  tag_117 = _RAND_117[19:0];
  _RAND_118 = {1{`RANDOM}};
  tag_118 = _RAND_118[19:0];
  _RAND_119 = {1{`RANDOM}};
  tag_119 = _RAND_119[19:0];
  _RAND_120 = {1{`RANDOM}};
  tag_120 = _RAND_120[19:0];
  _RAND_121 = {1{`RANDOM}};
  tag_121 = _RAND_121[19:0];
  _RAND_122 = {1{`RANDOM}};
  tag_122 = _RAND_122[19:0];
  _RAND_123 = {1{`RANDOM}};
  tag_123 = _RAND_123[19:0];
  _RAND_124 = {1{`RANDOM}};
  tag_124 = _RAND_124[19:0];
  _RAND_125 = {1{`RANDOM}};
  tag_125 = _RAND_125[19:0];
  _RAND_126 = {1{`RANDOM}};
  tag_126 = _RAND_126[19:0];
  _RAND_127 = {1{`RANDOM}};
  tag_127 = _RAND_127[19:0];
  _RAND_128 = {1{`RANDOM}};
  tag_128 = _RAND_128[19:0];
  _RAND_129 = {1{`RANDOM}};
  tag_129 = _RAND_129[19:0];
  _RAND_130 = {1{`RANDOM}};
  tag_130 = _RAND_130[19:0];
  _RAND_131 = {1{`RANDOM}};
  tag_131 = _RAND_131[19:0];
  _RAND_132 = {1{`RANDOM}};
  tag_132 = _RAND_132[19:0];
  _RAND_133 = {1{`RANDOM}};
  tag_133 = _RAND_133[19:0];
  _RAND_134 = {1{`RANDOM}};
  tag_134 = _RAND_134[19:0];
  _RAND_135 = {1{`RANDOM}};
  tag_135 = _RAND_135[19:0];
  _RAND_136 = {1{`RANDOM}};
  tag_136 = _RAND_136[19:0];
  _RAND_137 = {1{`RANDOM}};
  tag_137 = _RAND_137[19:0];
  _RAND_138 = {1{`RANDOM}};
  tag_138 = _RAND_138[19:0];
  _RAND_139 = {1{`RANDOM}};
  tag_139 = _RAND_139[19:0];
  _RAND_140 = {1{`RANDOM}};
  tag_140 = _RAND_140[19:0];
  _RAND_141 = {1{`RANDOM}};
  tag_141 = _RAND_141[19:0];
  _RAND_142 = {1{`RANDOM}};
  tag_142 = _RAND_142[19:0];
  _RAND_143 = {1{`RANDOM}};
  tag_143 = _RAND_143[19:0];
  _RAND_144 = {1{`RANDOM}};
  tag_144 = _RAND_144[19:0];
  _RAND_145 = {1{`RANDOM}};
  tag_145 = _RAND_145[19:0];
  _RAND_146 = {1{`RANDOM}};
  tag_146 = _RAND_146[19:0];
  _RAND_147 = {1{`RANDOM}};
  tag_147 = _RAND_147[19:0];
  _RAND_148 = {1{`RANDOM}};
  tag_148 = _RAND_148[19:0];
  _RAND_149 = {1{`RANDOM}};
  tag_149 = _RAND_149[19:0];
  _RAND_150 = {1{`RANDOM}};
  tag_150 = _RAND_150[19:0];
  _RAND_151 = {1{`RANDOM}};
  tag_151 = _RAND_151[19:0];
  _RAND_152 = {1{`RANDOM}};
  tag_152 = _RAND_152[19:0];
  _RAND_153 = {1{`RANDOM}};
  tag_153 = _RAND_153[19:0];
  _RAND_154 = {1{`RANDOM}};
  tag_154 = _RAND_154[19:0];
  _RAND_155 = {1{`RANDOM}};
  tag_155 = _RAND_155[19:0];
  _RAND_156 = {1{`RANDOM}};
  tag_156 = _RAND_156[19:0];
  _RAND_157 = {1{`RANDOM}};
  tag_157 = _RAND_157[19:0];
  _RAND_158 = {1{`RANDOM}};
  tag_158 = _RAND_158[19:0];
  _RAND_159 = {1{`RANDOM}};
  tag_159 = _RAND_159[19:0];
  _RAND_160 = {1{`RANDOM}};
  tag_160 = _RAND_160[19:0];
  _RAND_161 = {1{`RANDOM}};
  tag_161 = _RAND_161[19:0];
  _RAND_162 = {1{`RANDOM}};
  tag_162 = _RAND_162[19:0];
  _RAND_163 = {1{`RANDOM}};
  tag_163 = _RAND_163[19:0];
  _RAND_164 = {1{`RANDOM}};
  tag_164 = _RAND_164[19:0];
  _RAND_165 = {1{`RANDOM}};
  tag_165 = _RAND_165[19:0];
  _RAND_166 = {1{`RANDOM}};
  tag_166 = _RAND_166[19:0];
  _RAND_167 = {1{`RANDOM}};
  tag_167 = _RAND_167[19:0];
  _RAND_168 = {1{`RANDOM}};
  tag_168 = _RAND_168[19:0];
  _RAND_169 = {1{`RANDOM}};
  tag_169 = _RAND_169[19:0];
  _RAND_170 = {1{`RANDOM}};
  tag_170 = _RAND_170[19:0];
  _RAND_171 = {1{`RANDOM}};
  tag_171 = _RAND_171[19:0];
  _RAND_172 = {1{`RANDOM}};
  tag_172 = _RAND_172[19:0];
  _RAND_173 = {1{`RANDOM}};
  tag_173 = _RAND_173[19:0];
  _RAND_174 = {1{`RANDOM}};
  tag_174 = _RAND_174[19:0];
  _RAND_175 = {1{`RANDOM}};
  tag_175 = _RAND_175[19:0];
  _RAND_176 = {1{`RANDOM}};
  tag_176 = _RAND_176[19:0];
  _RAND_177 = {1{`RANDOM}};
  tag_177 = _RAND_177[19:0];
  _RAND_178 = {1{`RANDOM}};
  tag_178 = _RAND_178[19:0];
  _RAND_179 = {1{`RANDOM}};
  tag_179 = _RAND_179[19:0];
  _RAND_180 = {1{`RANDOM}};
  tag_180 = _RAND_180[19:0];
  _RAND_181 = {1{`RANDOM}};
  tag_181 = _RAND_181[19:0];
  _RAND_182 = {1{`RANDOM}};
  tag_182 = _RAND_182[19:0];
  _RAND_183 = {1{`RANDOM}};
  tag_183 = _RAND_183[19:0];
  _RAND_184 = {1{`RANDOM}};
  tag_184 = _RAND_184[19:0];
  _RAND_185 = {1{`RANDOM}};
  tag_185 = _RAND_185[19:0];
  _RAND_186 = {1{`RANDOM}};
  tag_186 = _RAND_186[19:0];
  _RAND_187 = {1{`RANDOM}};
  tag_187 = _RAND_187[19:0];
  _RAND_188 = {1{`RANDOM}};
  tag_188 = _RAND_188[19:0];
  _RAND_189 = {1{`RANDOM}};
  tag_189 = _RAND_189[19:0];
  _RAND_190 = {1{`RANDOM}};
  tag_190 = _RAND_190[19:0];
  _RAND_191 = {1{`RANDOM}};
  tag_191 = _RAND_191[19:0];
  _RAND_192 = {1{`RANDOM}};
  tag_192 = _RAND_192[19:0];
  _RAND_193 = {1{`RANDOM}};
  tag_193 = _RAND_193[19:0];
  _RAND_194 = {1{`RANDOM}};
  tag_194 = _RAND_194[19:0];
  _RAND_195 = {1{`RANDOM}};
  tag_195 = _RAND_195[19:0];
  _RAND_196 = {1{`RANDOM}};
  tag_196 = _RAND_196[19:0];
  _RAND_197 = {1{`RANDOM}};
  tag_197 = _RAND_197[19:0];
  _RAND_198 = {1{`RANDOM}};
  tag_198 = _RAND_198[19:0];
  _RAND_199 = {1{`RANDOM}};
  tag_199 = _RAND_199[19:0];
  _RAND_200 = {1{`RANDOM}};
  tag_200 = _RAND_200[19:0];
  _RAND_201 = {1{`RANDOM}};
  tag_201 = _RAND_201[19:0];
  _RAND_202 = {1{`RANDOM}};
  tag_202 = _RAND_202[19:0];
  _RAND_203 = {1{`RANDOM}};
  tag_203 = _RAND_203[19:0];
  _RAND_204 = {1{`RANDOM}};
  tag_204 = _RAND_204[19:0];
  _RAND_205 = {1{`RANDOM}};
  tag_205 = _RAND_205[19:0];
  _RAND_206 = {1{`RANDOM}};
  tag_206 = _RAND_206[19:0];
  _RAND_207 = {1{`RANDOM}};
  tag_207 = _RAND_207[19:0];
  _RAND_208 = {1{`RANDOM}};
  tag_208 = _RAND_208[19:0];
  _RAND_209 = {1{`RANDOM}};
  tag_209 = _RAND_209[19:0];
  _RAND_210 = {1{`RANDOM}};
  tag_210 = _RAND_210[19:0];
  _RAND_211 = {1{`RANDOM}};
  tag_211 = _RAND_211[19:0];
  _RAND_212 = {1{`RANDOM}};
  tag_212 = _RAND_212[19:0];
  _RAND_213 = {1{`RANDOM}};
  tag_213 = _RAND_213[19:0];
  _RAND_214 = {1{`RANDOM}};
  tag_214 = _RAND_214[19:0];
  _RAND_215 = {1{`RANDOM}};
  tag_215 = _RAND_215[19:0];
  _RAND_216 = {1{`RANDOM}};
  tag_216 = _RAND_216[19:0];
  _RAND_217 = {1{`RANDOM}};
  tag_217 = _RAND_217[19:0];
  _RAND_218 = {1{`RANDOM}};
  tag_218 = _RAND_218[19:0];
  _RAND_219 = {1{`RANDOM}};
  tag_219 = _RAND_219[19:0];
  _RAND_220 = {1{`RANDOM}};
  tag_220 = _RAND_220[19:0];
  _RAND_221 = {1{`RANDOM}};
  tag_221 = _RAND_221[19:0];
  _RAND_222 = {1{`RANDOM}};
  tag_222 = _RAND_222[19:0];
  _RAND_223 = {1{`RANDOM}};
  tag_223 = _RAND_223[19:0];
  _RAND_224 = {1{`RANDOM}};
  tag_224 = _RAND_224[19:0];
  _RAND_225 = {1{`RANDOM}};
  tag_225 = _RAND_225[19:0];
  _RAND_226 = {1{`RANDOM}};
  tag_226 = _RAND_226[19:0];
  _RAND_227 = {1{`RANDOM}};
  tag_227 = _RAND_227[19:0];
  _RAND_228 = {1{`RANDOM}};
  tag_228 = _RAND_228[19:0];
  _RAND_229 = {1{`RANDOM}};
  tag_229 = _RAND_229[19:0];
  _RAND_230 = {1{`RANDOM}};
  tag_230 = _RAND_230[19:0];
  _RAND_231 = {1{`RANDOM}};
  tag_231 = _RAND_231[19:0];
  _RAND_232 = {1{`RANDOM}};
  tag_232 = _RAND_232[19:0];
  _RAND_233 = {1{`RANDOM}};
  tag_233 = _RAND_233[19:0];
  _RAND_234 = {1{`RANDOM}};
  tag_234 = _RAND_234[19:0];
  _RAND_235 = {1{`RANDOM}};
  tag_235 = _RAND_235[19:0];
  _RAND_236 = {1{`RANDOM}};
  tag_236 = _RAND_236[19:0];
  _RAND_237 = {1{`RANDOM}};
  tag_237 = _RAND_237[19:0];
  _RAND_238 = {1{`RANDOM}};
  tag_238 = _RAND_238[19:0];
  _RAND_239 = {1{`RANDOM}};
  tag_239 = _RAND_239[19:0];
  _RAND_240 = {1{`RANDOM}};
  tag_240 = _RAND_240[19:0];
  _RAND_241 = {1{`RANDOM}};
  tag_241 = _RAND_241[19:0];
  _RAND_242 = {1{`RANDOM}};
  tag_242 = _RAND_242[19:0];
  _RAND_243 = {1{`RANDOM}};
  tag_243 = _RAND_243[19:0];
  _RAND_244 = {1{`RANDOM}};
  tag_244 = _RAND_244[19:0];
  _RAND_245 = {1{`RANDOM}};
  tag_245 = _RAND_245[19:0];
  _RAND_246 = {1{`RANDOM}};
  tag_246 = _RAND_246[19:0];
  _RAND_247 = {1{`RANDOM}};
  tag_247 = _RAND_247[19:0];
  _RAND_248 = {1{`RANDOM}};
  tag_248 = _RAND_248[19:0];
  _RAND_249 = {1{`RANDOM}};
  tag_249 = _RAND_249[19:0];
  _RAND_250 = {1{`RANDOM}};
  tag_250 = _RAND_250[19:0];
  _RAND_251 = {1{`RANDOM}};
  tag_251 = _RAND_251[19:0];
  _RAND_252 = {1{`RANDOM}};
  tag_252 = _RAND_252[19:0];
  _RAND_253 = {1{`RANDOM}};
  tag_253 = _RAND_253[19:0];
  _RAND_254 = {1{`RANDOM}};
  tag_254 = _RAND_254[19:0];
  _RAND_255 = {1{`RANDOM}};
  tag_255 = _RAND_255[19:0];
  _RAND_256 = {1{`RANDOM}};
  valid_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_3 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_4 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_5 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_6 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_7 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_8 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_9 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_10 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_11 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_12 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_13 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_14 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_15 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_16 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_17 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_18 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_19 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_20 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_21 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_22 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_23 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_24 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_25 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_26 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_27 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_28 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_29 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_30 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_31 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_32 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_33 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_34 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_35 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_36 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_37 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_38 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_39 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_40 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_41 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_42 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_43 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_44 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_45 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_46 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_47 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_48 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_49 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_50 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_51 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_52 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_53 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_54 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_55 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_56 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_57 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_58 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_59 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_60 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_61 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_62 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_63 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_64 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_65 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_66 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_67 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid_68 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid_69 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid_70 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid_71 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid_72 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid_73 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid_74 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid_75 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid_76 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid_77 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid_78 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid_79 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid_80 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid_81 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid_82 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid_83 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid_84 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid_85 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid_86 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid_87 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid_88 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid_89 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid_90 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid_91 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid_92 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid_93 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid_94 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid_95 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid_96 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid_97 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid_98 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid_99 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid_100 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid_101 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid_102 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid_103 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid_104 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid_105 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid_106 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid_107 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid_108 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid_109 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid_110 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid_111 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid_112 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid_113 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid_114 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid_115 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid_116 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid_117 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid_118 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid_119 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid_120 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid_121 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid_122 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid_123 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid_124 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid_125 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid_126 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid_127 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  valid_128 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  valid_129 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  valid_130 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  valid_131 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  valid_132 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  valid_133 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  valid_134 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  valid_135 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  valid_136 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  valid_137 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  valid_138 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  valid_139 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  valid_140 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  valid_141 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  valid_142 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  valid_143 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  valid_144 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  valid_145 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  valid_146 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  valid_147 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  valid_148 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  valid_149 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  valid_150 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  valid_151 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  valid_152 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  valid_153 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  valid_154 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  valid_155 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  valid_156 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  valid_157 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  valid_158 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  valid_159 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  valid_160 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  valid_161 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  valid_162 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  valid_163 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  valid_164 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  valid_165 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  valid_166 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  valid_167 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  valid_168 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  valid_169 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  valid_170 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  valid_171 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  valid_172 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  valid_173 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  valid_174 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  valid_175 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  valid_176 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  valid_177 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  valid_178 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  valid_179 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  valid_180 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  valid_181 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  valid_182 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  valid_183 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  valid_184 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  valid_185 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  valid_186 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  valid_187 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  valid_188 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  valid_189 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  valid_190 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  valid_191 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  valid_192 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  valid_193 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  valid_194 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  valid_195 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  valid_196 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  valid_197 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  valid_198 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  valid_199 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  valid_200 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  valid_201 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  valid_202 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  valid_203 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  valid_204 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  valid_205 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  valid_206 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  valid_207 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  valid_208 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  valid_209 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  valid_210 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  valid_211 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  valid_212 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  valid_213 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  valid_214 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  valid_215 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  valid_216 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  valid_217 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  valid_218 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  valid_219 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  valid_220 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  valid_221 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  valid_222 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  valid_223 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  valid_224 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  valid_225 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  valid_226 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  valid_227 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  valid_228 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  valid_229 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  valid_230 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  valid_231 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  valid_232 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  valid_233 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  valid_234 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  valid_235 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  valid_236 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  valid_237 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  valid_238 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  valid_239 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  valid_240 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  valid_241 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  valid_242 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  valid_243 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  valid_244 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  valid_245 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  valid_246 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  valid_247 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  valid_248 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  valid_249 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  valid_250 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  valid_251 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  valid_252 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  valid_253 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  valid_254 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  valid_255 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  dirty_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  dirty_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  dirty_2 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  dirty_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  dirty_4 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  dirty_5 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  dirty_6 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  dirty_7 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  dirty_8 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  dirty_9 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  dirty_10 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  dirty_11 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  dirty_12 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  dirty_13 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  dirty_14 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  dirty_15 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  dirty_16 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  dirty_17 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  dirty_18 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  dirty_19 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  dirty_20 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  dirty_21 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  dirty_22 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  dirty_23 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  dirty_24 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  dirty_25 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  dirty_26 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  dirty_27 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  dirty_28 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  dirty_29 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  dirty_30 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  dirty_31 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  dirty_32 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  dirty_33 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  dirty_34 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  dirty_35 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  dirty_36 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  dirty_37 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  dirty_38 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  dirty_39 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  dirty_40 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  dirty_41 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  dirty_42 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  dirty_43 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  dirty_44 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  dirty_45 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  dirty_46 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  dirty_47 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  dirty_48 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  dirty_49 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  dirty_50 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  dirty_51 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  dirty_52 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  dirty_53 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  dirty_54 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  dirty_55 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  dirty_56 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  dirty_57 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  dirty_58 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  dirty_59 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  dirty_60 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  dirty_61 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  dirty_62 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  dirty_63 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  dirty_64 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  dirty_65 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  dirty_66 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  dirty_67 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  dirty_68 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  dirty_69 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  dirty_70 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  dirty_71 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  dirty_72 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  dirty_73 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  dirty_74 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  dirty_75 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  dirty_76 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  dirty_77 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  dirty_78 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  dirty_79 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  dirty_80 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  dirty_81 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  dirty_82 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  dirty_83 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  dirty_84 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  dirty_85 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  dirty_86 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  dirty_87 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  dirty_88 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  dirty_89 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  dirty_90 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  dirty_91 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  dirty_92 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  dirty_93 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  dirty_94 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  dirty_95 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  dirty_96 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  dirty_97 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  dirty_98 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  dirty_99 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  dirty_100 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  dirty_101 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  dirty_102 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  dirty_103 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  dirty_104 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  dirty_105 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  dirty_106 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  dirty_107 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  dirty_108 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  dirty_109 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  dirty_110 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  dirty_111 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  dirty_112 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  dirty_113 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  dirty_114 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  dirty_115 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  dirty_116 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  dirty_117 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  dirty_118 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  dirty_119 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  dirty_120 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  dirty_121 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  dirty_122 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  dirty_123 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  dirty_124 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  dirty_125 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  dirty_126 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  dirty_127 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  dirty_128 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  dirty_129 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  dirty_130 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  dirty_131 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  dirty_132 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  dirty_133 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  dirty_134 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  dirty_135 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  dirty_136 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  dirty_137 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  dirty_138 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  dirty_139 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  dirty_140 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  dirty_141 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  dirty_142 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  dirty_143 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  dirty_144 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  dirty_145 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  dirty_146 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  dirty_147 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  dirty_148 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  dirty_149 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  dirty_150 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  dirty_151 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  dirty_152 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  dirty_153 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  dirty_154 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  dirty_155 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  dirty_156 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  dirty_157 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  dirty_158 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  dirty_159 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  dirty_160 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  dirty_161 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  dirty_162 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  dirty_163 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  dirty_164 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  dirty_165 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  dirty_166 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  dirty_167 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  dirty_168 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  dirty_169 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  dirty_170 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  dirty_171 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  dirty_172 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  dirty_173 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  dirty_174 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  dirty_175 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  dirty_176 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  dirty_177 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  dirty_178 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  dirty_179 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  dirty_180 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  dirty_181 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  dirty_182 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  dirty_183 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  dirty_184 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  dirty_185 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  dirty_186 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  dirty_187 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  dirty_188 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  dirty_189 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  dirty_190 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  dirty_191 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  dirty_192 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  dirty_193 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  dirty_194 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  dirty_195 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  dirty_196 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  dirty_197 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  dirty_198 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  dirty_199 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  dirty_200 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  dirty_201 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  dirty_202 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  dirty_203 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  dirty_204 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  dirty_205 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  dirty_206 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  dirty_207 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  dirty_208 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  dirty_209 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  dirty_210 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  dirty_211 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  dirty_212 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  dirty_213 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  dirty_214 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  dirty_215 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  dirty_216 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  dirty_217 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  dirty_218 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  dirty_219 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  dirty_220 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  dirty_221 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  dirty_222 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  dirty_223 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  dirty_224 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  dirty_225 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  dirty_226 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  dirty_227 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  dirty_228 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  dirty_229 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  dirty_230 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  dirty_231 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  dirty_232 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  dirty_233 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  dirty_234 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  dirty_235 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  dirty_236 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  dirty_237 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  dirty_238 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  dirty_239 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  dirty_240 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  dirty_241 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  dirty_242 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  dirty_243 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  dirty_244 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  dirty_245 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  dirty_246 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  dirty_247 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  dirty_248 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  dirty_249 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  dirty_250 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  dirty_251 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  dirty_252 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  dirty_253 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  dirty_254 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  dirty_255 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  offset_0 = _RAND_768[3:0];
  _RAND_769 = {1{`RANDOM}};
  offset_1 = _RAND_769[3:0];
  _RAND_770 = {1{`RANDOM}};
  offset_2 = _RAND_770[3:0];
  _RAND_771 = {1{`RANDOM}};
  offset_3 = _RAND_771[3:0];
  _RAND_772 = {1{`RANDOM}};
  offset_4 = _RAND_772[3:0];
  _RAND_773 = {1{`RANDOM}};
  offset_5 = _RAND_773[3:0];
  _RAND_774 = {1{`RANDOM}};
  offset_6 = _RAND_774[3:0];
  _RAND_775 = {1{`RANDOM}};
  offset_7 = _RAND_775[3:0];
  _RAND_776 = {1{`RANDOM}};
  offset_8 = _RAND_776[3:0];
  _RAND_777 = {1{`RANDOM}};
  offset_9 = _RAND_777[3:0];
  _RAND_778 = {1{`RANDOM}};
  offset_10 = _RAND_778[3:0];
  _RAND_779 = {1{`RANDOM}};
  offset_11 = _RAND_779[3:0];
  _RAND_780 = {1{`RANDOM}};
  offset_12 = _RAND_780[3:0];
  _RAND_781 = {1{`RANDOM}};
  offset_13 = _RAND_781[3:0];
  _RAND_782 = {1{`RANDOM}};
  offset_14 = _RAND_782[3:0];
  _RAND_783 = {1{`RANDOM}};
  offset_15 = _RAND_783[3:0];
  _RAND_784 = {1{`RANDOM}};
  offset_16 = _RAND_784[3:0];
  _RAND_785 = {1{`RANDOM}};
  offset_17 = _RAND_785[3:0];
  _RAND_786 = {1{`RANDOM}};
  offset_18 = _RAND_786[3:0];
  _RAND_787 = {1{`RANDOM}};
  offset_19 = _RAND_787[3:0];
  _RAND_788 = {1{`RANDOM}};
  offset_20 = _RAND_788[3:0];
  _RAND_789 = {1{`RANDOM}};
  offset_21 = _RAND_789[3:0];
  _RAND_790 = {1{`RANDOM}};
  offset_22 = _RAND_790[3:0];
  _RAND_791 = {1{`RANDOM}};
  offset_23 = _RAND_791[3:0];
  _RAND_792 = {1{`RANDOM}};
  offset_24 = _RAND_792[3:0];
  _RAND_793 = {1{`RANDOM}};
  offset_25 = _RAND_793[3:0];
  _RAND_794 = {1{`RANDOM}};
  offset_26 = _RAND_794[3:0];
  _RAND_795 = {1{`RANDOM}};
  offset_27 = _RAND_795[3:0];
  _RAND_796 = {1{`RANDOM}};
  offset_28 = _RAND_796[3:0];
  _RAND_797 = {1{`RANDOM}};
  offset_29 = _RAND_797[3:0];
  _RAND_798 = {1{`RANDOM}};
  offset_30 = _RAND_798[3:0];
  _RAND_799 = {1{`RANDOM}};
  offset_31 = _RAND_799[3:0];
  _RAND_800 = {1{`RANDOM}};
  offset_32 = _RAND_800[3:0];
  _RAND_801 = {1{`RANDOM}};
  offset_33 = _RAND_801[3:0];
  _RAND_802 = {1{`RANDOM}};
  offset_34 = _RAND_802[3:0];
  _RAND_803 = {1{`RANDOM}};
  offset_35 = _RAND_803[3:0];
  _RAND_804 = {1{`RANDOM}};
  offset_36 = _RAND_804[3:0];
  _RAND_805 = {1{`RANDOM}};
  offset_37 = _RAND_805[3:0];
  _RAND_806 = {1{`RANDOM}};
  offset_38 = _RAND_806[3:0];
  _RAND_807 = {1{`RANDOM}};
  offset_39 = _RAND_807[3:0];
  _RAND_808 = {1{`RANDOM}};
  offset_40 = _RAND_808[3:0];
  _RAND_809 = {1{`RANDOM}};
  offset_41 = _RAND_809[3:0];
  _RAND_810 = {1{`RANDOM}};
  offset_42 = _RAND_810[3:0];
  _RAND_811 = {1{`RANDOM}};
  offset_43 = _RAND_811[3:0];
  _RAND_812 = {1{`RANDOM}};
  offset_44 = _RAND_812[3:0];
  _RAND_813 = {1{`RANDOM}};
  offset_45 = _RAND_813[3:0];
  _RAND_814 = {1{`RANDOM}};
  offset_46 = _RAND_814[3:0];
  _RAND_815 = {1{`RANDOM}};
  offset_47 = _RAND_815[3:0];
  _RAND_816 = {1{`RANDOM}};
  offset_48 = _RAND_816[3:0];
  _RAND_817 = {1{`RANDOM}};
  offset_49 = _RAND_817[3:0];
  _RAND_818 = {1{`RANDOM}};
  offset_50 = _RAND_818[3:0];
  _RAND_819 = {1{`RANDOM}};
  offset_51 = _RAND_819[3:0];
  _RAND_820 = {1{`RANDOM}};
  offset_52 = _RAND_820[3:0];
  _RAND_821 = {1{`RANDOM}};
  offset_53 = _RAND_821[3:0];
  _RAND_822 = {1{`RANDOM}};
  offset_54 = _RAND_822[3:0];
  _RAND_823 = {1{`RANDOM}};
  offset_55 = _RAND_823[3:0];
  _RAND_824 = {1{`RANDOM}};
  offset_56 = _RAND_824[3:0];
  _RAND_825 = {1{`RANDOM}};
  offset_57 = _RAND_825[3:0];
  _RAND_826 = {1{`RANDOM}};
  offset_58 = _RAND_826[3:0];
  _RAND_827 = {1{`RANDOM}};
  offset_59 = _RAND_827[3:0];
  _RAND_828 = {1{`RANDOM}};
  offset_60 = _RAND_828[3:0];
  _RAND_829 = {1{`RANDOM}};
  offset_61 = _RAND_829[3:0];
  _RAND_830 = {1{`RANDOM}};
  offset_62 = _RAND_830[3:0];
  _RAND_831 = {1{`RANDOM}};
  offset_63 = _RAND_831[3:0];
  _RAND_832 = {1{`RANDOM}};
  offset_64 = _RAND_832[3:0];
  _RAND_833 = {1{`RANDOM}};
  offset_65 = _RAND_833[3:0];
  _RAND_834 = {1{`RANDOM}};
  offset_66 = _RAND_834[3:0];
  _RAND_835 = {1{`RANDOM}};
  offset_67 = _RAND_835[3:0];
  _RAND_836 = {1{`RANDOM}};
  offset_68 = _RAND_836[3:0];
  _RAND_837 = {1{`RANDOM}};
  offset_69 = _RAND_837[3:0];
  _RAND_838 = {1{`RANDOM}};
  offset_70 = _RAND_838[3:0];
  _RAND_839 = {1{`RANDOM}};
  offset_71 = _RAND_839[3:0];
  _RAND_840 = {1{`RANDOM}};
  offset_72 = _RAND_840[3:0];
  _RAND_841 = {1{`RANDOM}};
  offset_73 = _RAND_841[3:0];
  _RAND_842 = {1{`RANDOM}};
  offset_74 = _RAND_842[3:0];
  _RAND_843 = {1{`RANDOM}};
  offset_75 = _RAND_843[3:0];
  _RAND_844 = {1{`RANDOM}};
  offset_76 = _RAND_844[3:0];
  _RAND_845 = {1{`RANDOM}};
  offset_77 = _RAND_845[3:0];
  _RAND_846 = {1{`RANDOM}};
  offset_78 = _RAND_846[3:0];
  _RAND_847 = {1{`RANDOM}};
  offset_79 = _RAND_847[3:0];
  _RAND_848 = {1{`RANDOM}};
  offset_80 = _RAND_848[3:0];
  _RAND_849 = {1{`RANDOM}};
  offset_81 = _RAND_849[3:0];
  _RAND_850 = {1{`RANDOM}};
  offset_82 = _RAND_850[3:0];
  _RAND_851 = {1{`RANDOM}};
  offset_83 = _RAND_851[3:0];
  _RAND_852 = {1{`RANDOM}};
  offset_84 = _RAND_852[3:0];
  _RAND_853 = {1{`RANDOM}};
  offset_85 = _RAND_853[3:0];
  _RAND_854 = {1{`RANDOM}};
  offset_86 = _RAND_854[3:0];
  _RAND_855 = {1{`RANDOM}};
  offset_87 = _RAND_855[3:0];
  _RAND_856 = {1{`RANDOM}};
  offset_88 = _RAND_856[3:0];
  _RAND_857 = {1{`RANDOM}};
  offset_89 = _RAND_857[3:0];
  _RAND_858 = {1{`RANDOM}};
  offset_90 = _RAND_858[3:0];
  _RAND_859 = {1{`RANDOM}};
  offset_91 = _RAND_859[3:0];
  _RAND_860 = {1{`RANDOM}};
  offset_92 = _RAND_860[3:0];
  _RAND_861 = {1{`RANDOM}};
  offset_93 = _RAND_861[3:0];
  _RAND_862 = {1{`RANDOM}};
  offset_94 = _RAND_862[3:0];
  _RAND_863 = {1{`RANDOM}};
  offset_95 = _RAND_863[3:0];
  _RAND_864 = {1{`RANDOM}};
  offset_96 = _RAND_864[3:0];
  _RAND_865 = {1{`RANDOM}};
  offset_97 = _RAND_865[3:0];
  _RAND_866 = {1{`RANDOM}};
  offset_98 = _RAND_866[3:0];
  _RAND_867 = {1{`RANDOM}};
  offset_99 = _RAND_867[3:0];
  _RAND_868 = {1{`RANDOM}};
  offset_100 = _RAND_868[3:0];
  _RAND_869 = {1{`RANDOM}};
  offset_101 = _RAND_869[3:0];
  _RAND_870 = {1{`RANDOM}};
  offset_102 = _RAND_870[3:0];
  _RAND_871 = {1{`RANDOM}};
  offset_103 = _RAND_871[3:0];
  _RAND_872 = {1{`RANDOM}};
  offset_104 = _RAND_872[3:0];
  _RAND_873 = {1{`RANDOM}};
  offset_105 = _RAND_873[3:0];
  _RAND_874 = {1{`RANDOM}};
  offset_106 = _RAND_874[3:0];
  _RAND_875 = {1{`RANDOM}};
  offset_107 = _RAND_875[3:0];
  _RAND_876 = {1{`RANDOM}};
  offset_108 = _RAND_876[3:0];
  _RAND_877 = {1{`RANDOM}};
  offset_109 = _RAND_877[3:0];
  _RAND_878 = {1{`RANDOM}};
  offset_110 = _RAND_878[3:0];
  _RAND_879 = {1{`RANDOM}};
  offset_111 = _RAND_879[3:0];
  _RAND_880 = {1{`RANDOM}};
  offset_112 = _RAND_880[3:0];
  _RAND_881 = {1{`RANDOM}};
  offset_113 = _RAND_881[3:0];
  _RAND_882 = {1{`RANDOM}};
  offset_114 = _RAND_882[3:0];
  _RAND_883 = {1{`RANDOM}};
  offset_115 = _RAND_883[3:0];
  _RAND_884 = {1{`RANDOM}};
  offset_116 = _RAND_884[3:0];
  _RAND_885 = {1{`RANDOM}};
  offset_117 = _RAND_885[3:0];
  _RAND_886 = {1{`RANDOM}};
  offset_118 = _RAND_886[3:0];
  _RAND_887 = {1{`RANDOM}};
  offset_119 = _RAND_887[3:0];
  _RAND_888 = {1{`RANDOM}};
  offset_120 = _RAND_888[3:0];
  _RAND_889 = {1{`RANDOM}};
  offset_121 = _RAND_889[3:0];
  _RAND_890 = {1{`RANDOM}};
  offset_122 = _RAND_890[3:0];
  _RAND_891 = {1{`RANDOM}};
  offset_123 = _RAND_891[3:0];
  _RAND_892 = {1{`RANDOM}};
  offset_124 = _RAND_892[3:0];
  _RAND_893 = {1{`RANDOM}};
  offset_125 = _RAND_893[3:0];
  _RAND_894 = {1{`RANDOM}};
  offset_126 = _RAND_894[3:0];
  _RAND_895 = {1{`RANDOM}};
  offset_127 = _RAND_895[3:0];
  _RAND_896 = {1{`RANDOM}};
  offset_128 = _RAND_896[3:0];
  _RAND_897 = {1{`RANDOM}};
  offset_129 = _RAND_897[3:0];
  _RAND_898 = {1{`RANDOM}};
  offset_130 = _RAND_898[3:0];
  _RAND_899 = {1{`RANDOM}};
  offset_131 = _RAND_899[3:0];
  _RAND_900 = {1{`RANDOM}};
  offset_132 = _RAND_900[3:0];
  _RAND_901 = {1{`RANDOM}};
  offset_133 = _RAND_901[3:0];
  _RAND_902 = {1{`RANDOM}};
  offset_134 = _RAND_902[3:0];
  _RAND_903 = {1{`RANDOM}};
  offset_135 = _RAND_903[3:0];
  _RAND_904 = {1{`RANDOM}};
  offset_136 = _RAND_904[3:0];
  _RAND_905 = {1{`RANDOM}};
  offset_137 = _RAND_905[3:0];
  _RAND_906 = {1{`RANDOM}};
  offset_138 = _RAND_906[3:0];
  _RAND_907 = {1{`RANDOM}};
  offset_139 = _RAND_907[3:0];
  _RAND_908 = {1{`RANDOM}};
  offset_140 = _RAND_908[3:0];
  _RAND_909 = {1{`RANDOM}};
  offset_141 = _RAND_909[3:0];
  _RAND_910 = {1{`RANDOM}};
  offset_142 = _RAND_910[3:0];
  _RAND_911 = {1{`RANDOM}};
  offset_143 = _RAND_911[3:0];
  _RAND_912 = {1{`RANDOM}};
  offset_144 = _RAND_912[3:0];
  _RAND_913 = {1{`RANDOM}};
  offset_145 = _RAND_913[3:0];
  _RAND_914 = {1{`RANDOM}};
  offset_146 = _RAND_914[3:0];
  _RAND_915 = {1{`RANDOM}};
  offset_147 = _RAND_915[3:0];
  _RAND_916 = {1{`RANDOM}};
  offset_148 = _RAND_916[3:0];
  _RAND_917 = {1{`RANDOM}};
  offset_149 = _RAND_917[3:0];
  _RAND_918 = {1{`RANDOM}};
  offset_150 = _RAND_918[3:0];
  _RAND_919 = {1{`RANDOM}};
  offset_151 = _RAND_919[3:0];
  _RAND_920 = {1{`RANDOM}};
  offset_152 = _RAND_920[3:0];
  _RAND_921 = {1{`RANDOM}};
  offset_153 = _RAND_921[3:0];
  _RAND_922 = {1{`RANDOM}};
  offset_154 = _RAND_922[3:0];
  _RAND_923 = {1{`RANDOM}};
  offset_155 = _RAND_923[3:0];
  _RAND_924 = {1{`RANDOM}};
  offset_156 = _RAND_924[3:0];
  _RAND_925 = {1{`RANDOM}};
  offset_157 = _RAND_925[3:0];
  _RAND_926 = {1{`RANDOM}};
  offset_158 = _RAND_926[3:0];
  _RAND_927 = {1{`RANDOM}};
  offset_159 = _RAND_927[3:0];
  _RAND_928 = {1{`RANDOM}};
  offset_160 = _RAND_928[3:0];
  _RAND_929 = {1{`RANDOM}};
  offset_161 = _RAND_929[3:0];
  _RAND_930 = {1{`RANDOM}};
  offset_162 = _RAND_930[3:0];
  _RAND_931 = {1{`RANDOM}};
  offset_163 = _RAND_931[3:0];
  _RAND_932 = {1{`RANDOM}};
  offset_164 = _RAND_932[3:0];
  _RAND_933 = {1{`RANDOM}};
  offset_165 = _RAND_933[3:0];
  _RAND_934 = {1{`RANDOM}};
  offset_166 = _RAND_934[3:0];
  _RAND_935 = {1{`RANDOM}};
  offset_167 = _RAND_935[3:0];
  _RAND_936 = {1{`RANDOM}};
  offset_168 = _RAND_936[3:0];
  _RAND_937 = {1{`RANDOM}};
  offset_169 = _RAND_937[3:0];
  _RAND_938 = {1{`RANDOM}};
  offset_170 = _RAND_938[3:0];
  _RAND_939 = {1{`RANDOM}};
  offset_171 = _RAND_939[3:0];
  _RAND_940 = {1{`RANDOM}};
  offset_172 = _RAND_940[3:0];
  _RAND_941 = {1{`RANDOM}};
  offset_173 = _RAND_941[3:0];
  _RAND_942 = {1{`RANDOM}};
  offset_174 = _RAND_942[3:0];
  _RAND_943 = {1{`RANDOM}};
  offset_175 = _RAND_943[3:0];
  _RAND_944 = {1{`RANDOM}};
  offset_176 = _RAND_944[3:0];
  _RAND_945 = {1{`RANDOM}};
  offset_177 = _RAND_945[3:0];
  _RAND_946 = {1{`RANDOM}};
  offset_178 = _RAND_946[3:0];
  _RAND_947 = {1{`RANDOM}};
  offset_179 = _RAND_947[3:0];
  _RAND_948 = {1{`RANDOM}};
  offset_180 = _RAND_948[3:0];
  _RAND_949 = {1{`RANDOM}};
  offset_181 = _RAND_949[3:0];
  _RAND_950 = {1{`RANDOM}};
  offset_182 = _RAND_950[3:0];
  _RAND_951 = {1{`RANDOM}};
  offset_183 = _RAND_951[3:0];
  _RAND_952 = {1{`RANDOM}};
  offset_184 = _RAND_952[3:0];
  _RAND_953 = {1{`RANDOM}};
  offset_185 = _RAND_953[3:0];
  _RAND_954 = {1{`RANDOM}};
  offset_186 = _RAND_954[3:0];
  _RAND_955 = {1{`RANDOM}};
  offset_187 = _RAND_955[3:0];
  _RAND_956 = {1{`RANDOM}};
  offset_188 = _RAND_956[3:0];
  _RAND_957 = {1{`RANDOM}};
  offset_189 = _RAND_957[3:0];
  _RAND_958 = {1{`RANDOM}};
  offset_190 = _RAND_958[3:0];
  _RAND_959 = {1{`RANDOM}};
  offset_191 = _RAND_959[3:0];
  _RAND_960 = {1{`RANDOM}};
  offset_192 = _RAND_960[3:0];
  _RAND_961 = {1{`RANDOM}};
  offset_193 = _RAND_961[3:0];
  _RAND_962 = {1{`RANDOM}};
  offset_194 = _RAND_962[3:0];
  _RAND_963 = {1{`RANDOM}};
  offset_195 = _RAND_963[3:0];
  _RAND_964 = {1{`RANDOM}};
  offset_196 = _RAND_964[3:0];
  _RAND_965 = {1{`RANDOM}};
  offset_197 = _RAND_965[3:0];
  _RAND_966 = {1{`RANDOM}};
  offset_198 = _RAND_966[3:0];
  _RAND_967 = {1{`RANDOM}};
  offset_199 = _RAND_967[3:0];
  _RAND_968 = {1{`RANDOM}};
  offset_200 = _RAND_968[3:0];
  _RAND_969 = {1{`RANDOM}};
  offset_201 = _RAND_969[3:0];
  _RAND_970 = {1{`RANDOM}};
  offset_202 = _RAND_970[3:0];
  _RAND_971 = {1{`RANDOM}};
  offset_203 = _RAND_971[3:0];
  _RAND_972 = {1{`RANDOM}};
  offset_204 = _RAND_972[3:0];
  _RAND_973 = {1{`RANDOM}};
  offset_205 = _RAND_973[3:0];
  _RAND_974 = {1{`RANDOM}};
  offset_206 = _RAND_974[3:0];
  _RAND_975 = {1{`RANDOM}};
  offset_207 = _RAND_975[3:0];
  _RAND_976 = {1{`RANDOM}};
  offset_208 = _RAND_976[3:0];
  _RAND_977 = {1{`RANDOM}};
  offset_209 = _RAND_977[3:0];
  _RAND_978 = {1{`RANDOM}};
  offset_210 = _RAND_978[3:0];
  _RAND_979 = {1{`RANDOM}};
  offset_211 = _RAND_979[3:0];
  _RAND_980 = {1{`RANDOM}};
  offset_212 = _RAND_980[3:0];
  _RAND_981 = {1{`RANDOM}};
  offset_213 = _RAND_981[3:0];
  _RAND_982 = {1{`RANDOM}};
  offset_214 = _RAND_982[3:0];
  _RAND_983 = {1{`RANDOM}};
  offset_215 = _RAND_983[3:0];
  _RAND_984 = {1{`RANDOM}};
  offset_216 = _RAND_984[3:0];
  _RAND_985 = {1{`RANDOM}};
  offset_217 = _RAND_985[3:0];
  _RAND_986 = {1{`RANDOM}};
  offset_218 = _RAND_986[3:0];
  _RAND_987 = {1{`RANDOM}};
  offset_219 = _RAND_987[3:0];
  _RAND_988 = {1{`RANDOM}};
  offset_220 = _RAND_988[3:0];
  _RAND_989 = {1{`RANDOM}};
  offset_221 = _RAND_989[3:0];
  _RAND_990 = {1{`RANDOM}};
  offset_222 = _RAND_990[3:0];
  _RAND_991 = {1{`RANDOM}};
  offset_223 = _RAND_991[3:0];
  _RAND_992 = {1{`RANDOM}};
  offset_224 = _RAND_992[3:0];
  _RAND_993 = {1{`RANDOM}};
  offset_225 = _RAND_993[3:0];
  _RAND_994 = {1{`RANDOM}};
  offset_226 = _RAND_994[3:0];
  _RAND_995 = {1{`RANDOM}};
  offset_227 = _RAND_995[3:0];
  _RAND_996 = {1{`RANDOM}};
  offset_228 = _RAND_996[3:0];
  _RAND_997 = {1{`RANDOM}};
  offset_229 = _RAND_997[3:0];
  _RAND_998 = {1{`RANDOM}};
  offset_230 = _RAND_998[3:0];
  _RAND_999 = {1{`RANDOM}};
  offset_231 = _RAND_999[3:0];
  _RAND_1000 = {1{`RANDOM}};
  offset_232 = _RAND_1000[3:0];
  _RAND_1001 = {1{`RANDOM}};
  offset_233 = _RAND_1001[3:0];
  _RAND_1002 = {1{`RANDOM}};
  offset_234 = _RAND_1002[3:0];
  _RAND_1003 = {1{`RANDOM}};
  offset_235 = _RAND_1003[3:0];
  _RAND_1004 = {1{`RANDOM}};
  offset_236 = _RAND_1004[3:0];
  _RAND_1005 = {1{`RANDOM}};
  offset_237 = _RAND_1005[3:0];
  _RAND_1006 = {1{`RANDOM}};
  offset_238 = _RAND_1006[3:0];
  _RAND_1007 = {1{`RANDOM}};
  offset_239 = _RAND_1007[3:0];
  _RAND_1008 = {1{`RANDOM}};
  offset_240 = _RAND_1008[3:0];
  _RAND_1009 = {1{`RANDOM}};
  offset_241 = _RAND_1009[3:0];
  _RAND_1010 = {1{`RANDOM}};
  offset_242 = _RAND_1010[3:0];
  _RAND_1011 = {1{`RANDOM}};
  offset_243 = _RAND_1011[3:0];
  _RAND_1012 = {1{`RANDOM}};
  offset_244 = _RAND_1012[3:0];
  _RAND_1013 = {1{`RANDOM}};
  offset_245 = _RAND_1013[3:0];
  _RAND_1014 = {1{`RANDOM}};
  offset_246 = _RAND_1014[3:0];
  _RAND_1015 = {1{`RANDOM}};
  offset_247 = _RAND_1015[3:0];
  _RAND_1016 = {1{`RANDOM}};
  offset_248 = _RAND_1016[3:0];
  _RAND_1017 = {1{`RANDOM}};
  offset_249 = _RAND_1017[3:0];
  _RAND_1018 = {1{`RANDOM}};
  offset_250 = _RAND_1018[3:0];
  _RAND_1019 = {1{`RANDOM}};
  offset_251 = _RAND_1019[3:0];
  _RAND_1020 = {1{`RANDOM}};
  offset_252 = _RAND_1020[3:0];
  _RAND_1021 = {1{`RANDOM}};
  offset_253 = _RAND_1021[3:0];
  _RAND_1022 = {1{`RANDOM}};
  offset_254 = _RAND_1022[3:0];
  _RAND_1023 = {1{`RANDOM}};
  offset_255 = _RAND_1023[3:0];
  _RAND_1024 = {1{`RANDOM}};
  state = _RAND_1024[2:0];
  _RAND_1025 = {1{`RANDOM}};
  data_ready = _RAND_1025[0:0];
  _RAND_1026 = {1{`RANDOM}};
  cache_fill = _RAND_1026[0:0];
  _RAND_1027 = {1{`RANDOM}};
  cache_wen = _RAND_1027[0:0];
  _RAND_1028 = {4{`RANDOM}};
  cache_wdata = _RAND_1028[127:0];
  _RAND_1029 = {4{`RANDOM}};
  cache_strb = _RAND_1029[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AxiLite2Axi(
  input          clock,
  input          reset,
  input          io_out_aw_ready,
  output         io_out_aw_valid,
  output [31:0]  io_out_aw_bits_addr,
  input          io_out_w_ready,
  output         io_out_w_valid,
  output [63:0]  io_out_w_bits_data,
  output [7:0]   io_out_w_bits_strb,
  output         io_out_w_bits_last,
  output         io_out_b_ready,
  input          io_out_b_valid,
  input          io_out_ar_ready,
  output         io_out_ar_valid,
  output [31:0]  io_out_ar_bits_addr,
  output         io_out_r_ready,
  input          io_out_r_valid,
  input  [63:0]  io_out_r_bits_data,
  input          io_out_r_bits_last,
  input          io_imem_inst_valid,
  output         io_imem_inst_ready,
  input  [31:0]  io_imem_inst_addr,
  output [127:0] io_imem_inst_read,
  input          io_dmem_data_valid,
  output         io_dmem_data_ready,
  input          io_dmem_data_req,
  input  [31:0]  io_dmem_data_addr,
  input  [7:0]   io_dmem_data_strb,
  output [127:0] io_dmem_data_read,
  input  [127:0] io_dmem_data_write
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  data_ren = io_dmem_data_valid & ~io_dmem_data_req; // @[AXI.scala 123:30]
  wire  data_wen = io_dmem_data_valid & io_dmem_data_req; // @[AXI.scala 124:30]
  wire  aw_hs = io_out_aw_ready & io_out_aw_valid; // @[AXI.scala 126:33]
  wire  w_hs = io_out_w_ready & io_out_w_valid; // @[AXI.scala 127:33]
  wire  b_hs = io_out_b_ready & io_out_b_valid; // @[AXI.scala 128:33]
  wire  ar_hs = io_out_ar_ready & io_out_ar_valid; // @[AXI.scala 129:33]
  wire  r_hs = io_out_r_ready & io_out_r_valid; // @[AXI.scala 130:33]
  wire  w_done = w_hs & io_out_w_bits_last; // @[AXI.scala 132:25]
  wire  r_done = r_hs & io_out_r_bits_last; // @[AXI.scala 133:25]
  reg [2:0] r_state; // @[AXI.scala 136:24]
  reg [2:0] w_state; // @[AXI.scala 139:24]
  wire  _T = 3'h0 == r_state; // @[Conditional.scala 37:30]
  wire  _T_1 = 3'h1 == r_state; // @[Conditional.scala 37:30]
  wire  _T_2 = 3'h2 == r_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_3 = r_done ? 3'h3 : r_state; // @[AXI.scala 156:21 AXI.scala 157:17 AXI.scala 136:24]
  wire  _T_3 = 3'h3 == r_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_4 = data_ren ? 3'h4 : 3'h0; // @[AXI.scala 161:23 AXI.scala 162:17 AXI.scala 165:17]
  wire  _T_4 = 3'h4 == r_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_5 = ar_hs ? 3'h5 : r_state; // @[AXI.scala 169:20 AXI.scala 170:17 AXI.scala 136:24]
  wire  _T_5 = 3'h5 == r_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_6 = r_done ? 3'h6 : r_state; // @[AXI.scala 174:21 AXI.scala 175:17 AXI.scala 136:24]
  wire  _T_6 = 3'h6 == r_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_7 = _T_6 ? 3'h0 : r_state; // @[Conditional.scala 39:67 AXI.scala 179:15 AXI.scala 136:24]
  wire [2:0] _GEN_8 = _T_5 ? _GEN_6 : _GEN_7; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_9 = _T_4 ? _GEN_5 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_3 ? _GEN_4 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _T_7 = 3'h0 == w_state; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h1 == w_state; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h2 == w_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_16 = w_done ? 3'h3 : w_state; // @[AXI.scala 195:21 AXI.scala 196:17 AXI.scala 139:24]
  wire  _T_10 = 3'h3 == w_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_17 = b_hs ? 3'h4 : w_state; // @[AXI.scala 200:19 AXI.scala 201:17 AXI.scala 139:24]
  wire  _T_11 = 3'h4 == w_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_18 = _T_11 ? 3'h0 : w_state; // @[Conditional.scala 39:67 AXI.scala 205:15 AXI.scala 139:24]
  wire [2:0] _GEN_19 = _T_10 ? _GEN_17 : _GEN_18; // @[Conditional.scala 39:67]
  reg  data_ok; // @[AXI.scala 209:24]
  wire  _T_12 = w_state == 3'h4; // @[AXI.scala 210:29]
  wire  _GEN_23 = ~data_wen ? 1'h0 : data_ok; // @[AXI.scala 213:25 AXI.scala 214:13 AXI.scala 209:24]
  wire  _GEN_24 = data_wen & w_state == 3'h4 | _GEN_23; // @[AXI.scala 210:46 AXI.scala 211:13]
  wire  _axi_addr_T = r_state == 3'h1; // @[AXI.scala 217:31]
  wire [31:0] _axi_addr_T_1 = io_imem_inst_addr & 32'hfffffff0; // @[AXI.scala 217:62]
  wire  _axi_addr_T_2 = r_state == 3'h4; // @[AXI.scala 218:31]
  wire [31:0] _axi_addr_T_3 = io_dmem_data_addr & 32'hfffffff0; // @[AXI.scala 218:62]
  wire [31:0] _axi_addr_T_4 = r_state == 3'h4 ? _axi_addr_T_3 : 32'h0; // @[AXI.scala 218:22]
  wire [27:0] axi_waddr_hi = io_dmem_data_addr[31:4]; // @[AXI.scala 219:49]
  wire [31:0] _axi_waddr_T = {axi_waddr_hi,4'h8}; // @[Cat.scala 30:58]
  reg [63:0] inst_read_h; // @[AXI.scala 265:28]
  reg [63:0] inst_read_l; // @[AXI.scala 266:28]
  reg [63:0] data_read_h; // @[AXI.scala 267:28]
  reg [63:0] data_read_l; // @[AXI.scala 268:28]
  assign io_out_aw_valid = w_state == 3'h1; // @[AXI.scala 238:34]
  assign io_out_aw_bits_addr = data_ok ? _axi_waddr_T : _axi_addr_T_3; // @[AXI.scala 219:22]
  assign io_out_w_valid = w_state == 3'h2; // @[AXI.scala 251:34]
  assign io_out_w_bits_data = data_ok ? io_dmem_data_write[127:64] : io_dmem_data_write[63:0]; // @[AXI.scala 252:29]
  assign io_out_w_bits_strb = io_dmem_data_strb; // @[AXI.scala 253:23]
  assign io_out_w_bits_last = 1'h1; // @[AXI.scala 254:23]
  assign io_out_b_ready = 1'h1; // @[AXI.scala 256:23]
  assign io_out_ar_valid = _axi_addr_T | _axi_addr_T_2; // @[AXI.scala 222:50]
  assign io_out_ar_bits_addr = r_state == 3'h1 ? _axi_addr_T_1 : _axi_addr_T_4; // @[AXI.scala 217:22]
  assign io_out_r_ready = 1'h1; // @[AXI.scala 235:23]
  assign io_imem_inst_ready = r_state == 3'h3; // @[AXI.scala 262:29]
  assign io_imem_inst_read = {inst_read_h,inst_read_l}; // @[Cat.scala 30:58]
  assign io_dmem_data_ready = r_state == 3'h6 | _T_12 & data_ok; // @[AXI.scala 263:45]
  assign io_dmem_data_read = {data_read_h,data_read_l}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if (reset) begin // @[AXI.scala 136:24]
      r_state <= 3'h0; // @[AXI.scala 136:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_imem_inst_valid) begin // @[AXI.scala 143:23]
        r_state <= 3'h1; // @[AXI.scala 144:17]
      end else if (data_ren) begin // @[AXI.scala 146:28]
        r_state <= 3'h4; // @[AXI.scala 147:17]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (ar_hs) begin // @[AXI.scala 151:20]
        r_state <= 3'h2; // @[AXI.scala 152:17]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      r_state <= _GEN_3;
    end else begin
      r_state <= _GEN_10;
    end
    if (reset) begin // @[AXI.scala 139:24]
      w_state <= 3'h0; // @[AXI.scala 139:24]
    end else if (_T_7) begin // @[Conditional.scala 40:58]
      if (data_wen) begin // @[AXI.scala 185:23]
        w_state <= 3'h1; // @[AXI.scala 186:17]
      end
    end else if (_T_8) begin // @[Conditional.scala 39:67]
      if (aw_hs) begin // @[AXI.scala 190:20]
        w_state <= 3'h2; // @[AXI.scala 191:17]
      end
    end else if (_T_9) begin // @[Conditional.scala 39:67]
      w_state <= _GEN_16;
    end else begin
      w_state <= _GEN_19;
    end
    if (reset) begin // @[AXI.scala 209:24]
      data_ok <= 1'h0; // @[AXI.scala 209:24]
    end else begin
      data_ok <= _GEN_24;
    end
    if (reset) begin // @[AXI.scala 265:28]
      inst_read_h <= 64'h0; // @[AXI.scala 265:28]
    end else if (r_hs) begin // @[AXI.scala 270:15]
      if (io_out_r_bits_last) begin // @[AXI.scala 271:28]
        inst_read_h <= io_out_r_bits_data; // @[AXI.scala 272:19]
      end
    end
    if (reset) begin // @[AXI.scala 266:28]
      inst_read_l <= 64'h0; // @[AXI.scala 266:28]
    end else if (r_hs) begin // @[AXI.scala 270:15]
      if (!(io_out_r_bits_last)) begin // @[AXI.scala 271:28]
        inst_read_l <= io_out_r_bits_data; // @[AXI.scala 276:19]
      end
    end
    if (reset) begin // @[AXI.scala 267:28]
      data_read_h <= 64'h0; // @[AXI.scala 267:28]
    end else if (r_hs) begin // @[AXI.scala 270:15]
      if (io_out_r_bits_last) begin // @[AXI.scala 271:28]
        data_read_h <= io_out_r_bits_data; // @[AXI.scala 273:19]
      end
    end
    if (reset) begin // @[AXI.scala 268:28]
      data_read_l <= 64'h0; // @[AXI.scala 268:28]
    end else if (r_hs) begin // @[AXI.scala 270:15]
      if (!(io_out_r_bits_last)) begin // @[AXI.scala 271:28]
        data_read_l <= io_out_r_bits_data; // @[AXI.scala 277:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  w_state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  data_ok = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  inst_read_h = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  inst_read_l = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  data_read_h = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  data_read_l = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimTop(
  input         clock,
  input         reset,
  input  [63:0] io_logCtrl_log_begin,
  input  [63:0] io_logCtrl_log_end,
  input  [63:0] io_logCtrl_log_level,
  input         io_perfInfo_clean,
  input         io_perfInfo_dump,
  output        io_uart_out_valid,
  output [7:0]  io_uart_out_ch,
  output        io_uart_in_valid,
  input  [7:0]  io_uart_in_ch,
  input         io_memAXI_0_aw_ready,
  output        io_memAXI_0_aw_valid,
  output [31:0] io_memAXI_0_aw_bits_addr,
  output [2:0]  io_memAXI_0_aw_bits_prot,
  output [3:0]  io_memAXI_0_aw_bits_id,
  output        io_memAXI_0_aw_bits_user,
  output [7:0]  io_memAXI_0_aw_bits_len,
  output [2:0]  io_memAXI_0_aw_bits_size,
  output [1:0]  io_memAXI_0_aw_bits_burst,
  output        io_memAXI_0_aw_bits_lock,
  output [3:0]  io_memAXI_0_aw_bits_cache,
  output [3:0]  io_memAXI_0_aw_bits_qos,
  input         io_memAXI_0_w_ready,
  output        io_memAXI_0_w_valid,
  output [63:0] io_memAXI_0_w_bits_data,
  output [7:0]  io_memAXI_0_w_bits_strb,
  output        io_memAXI_0_w_bits_last,
  output        io_memAXI_0_b_ready,
  input         io_memAXI_0_b_valid,
  input  [1:0]  io_memAXI_0_b_bits_resp,
  input  [3:0]  io_memAXI_0_b_bits_id,
  input         io_memAXI_0_b_bits_user,
  input         io_memAXI_0_ar_ready,
  output        io_memAXI_0_ar_valid,
  output [31:0] io_memAXI_0_ar_bits_addr,
  output [2:0]  io_memAXI_0_ar_bits_prot,
  output [3:0]  io_memAXI_0_ar_bits_id,
  output        io_memAXI_0_ar_bits_user,
  output [7:0]  io_memAXI_0_ar_bits_len,
  output [2:0]  io_memAXI_0_ar_bits_size,
  output [1:0]  io_memAXI_0_ar_bits_burst,
  output        io_memAXI_0_ar_bits_lock,
  output [3:0]  io_memAXI_0_ar_bits_cache,
  output [3:0]  io_memAXI_0_ar_bits_qos,
  output        io_memAXI_0_r_ready,
  input         io_memAXI_0_r_valid,
  input  [1:0]  io_memAXI_0_r_bits_resp,
  input  [63:0] io_memAXI_0_r_bits_data,
  input  [3:0]  io_memAXI_0_r_bits_id,
  input         io_memAXI_0_r_bits_user,
  input         io_memAXI_0_r_bits_last
);
  wire  core_clock; // @[SimTop.scala 15:20]
  wire  core_reset; // @[SimTop.scala 15:20]
  wire  core_io_imem_inst_valid; // @[SimTop.scala 15:20]
  wire  core_io_imem_inst_ready; // @[SimTop.scala 15:20]
  wire [31:0] core_io_imem_inst_addr; // @[SimTop.scala 15:20]
  wire [31:0] core_io_imem_inst_read; // @[SimTop.scala 15:20]
  wire  core_io_dmem_data_valid; // @[SimTop.scala 15:20]
  wire  core_io_dmem_data_ready; // @[SimTop.scala 15:20]
  wire  core_io_dmem_data_req; // @[SimTop.scala 15:20]
  wire [31:0] core_io_dmem_data_addr; // @[SimTop.scala 15:20]
  wire [1:0] core_io_dmem_data_size; // @[SimTop.scala 15:20]
  wire [7:0] core_io_dmem_data_strb; // @[SimTop.scala 15:20]
  wire [63:0] core_io_dmem_data_read; // @[SimTop.scala 15:20]
  wire [63:0] core_io_dmem_data_write; // @[SimTop.scala 15:20]
  wire  icache_clock; // @[SimTop.scala 16:22]
  wire  icache_reset; // @[SimTop.scala 16:22]
  wire  icache_io_imem_inst_valid; // @[SimTop.scala 16:22]
  wire  icache_io_imem_inst_ready; // @[SimTop.scala 16:22]
  wire [31:0] icache_io_imem_inst_addr; // @[SimTop.scala 16:22]
  wire [31:0] icache_io_imem_inst_read; // @[SimTop.scala 16:22]
  wire  icache_io_out_inst_valid; // @[SimTop.scala 16:22]
  wire  icache_io_out_inst_ready; // @[SimTop.scala 16:22]
  wire [31:0] icache_io_out_inst_addr; // @[SimTop.scala 16:22]
  wire [127:0] icache_io_out_inst_read; // @[SimTop.scala 16:22]
  wire  dcache_clock; // @[SimTop.scala 17:22]
  wire  dcache_reset; // @[SimTop.scala 17:22]
  wire  dcache_io_dmem_data_valid; // @[SimTop.scala 17:22]
  wire  dcache_io_dmem_data_ready; // @[SimTop.scala 17:22]
  wire  dcache_io_dmem_data_req; // @[SimTop.scala 17:22]
  wire [31:0] dcache_io_dmem_data_addr; // @[SimTop.scala 17:22]
  wire [1:0] dcache_io_dmem_data_size; // @[SimTop.scala 17:22]
  wire [7:0] dcache_io_dmem_data_strb; // @[SimTop.scala 17:22]
  wire [63:0] dcache_io_dmem_data_read; // @[SimTop.scala 17:22]
  wire [63:0] dcache_io_dmem_data_write; // @[SimTop.scala 17:22]
  wire  dcache_io_out_data_valid; // @[SimTop.scala 17:22]
  wire  dcache_io_out_data_ready; // @[SimTop.scala 17:22]
  wire  dcache_io_out_data_req; // @[SimTop.scala 17:22]
  wire [31:0] dcache_io_out_data_addr; // @[SimTop.scala 17:22]
  wire [7:0] dcache_io_out_data_strb; // @[SimTop.scala 17:22]
  wire [127:0] dcache_io_out_data_read; // @[SimTop.scala 17:22]
  wire [127:0] dcache_io_out_data_write; // @[SimTop.scala 17:22]
  wire  top_clock; // @[SimTop.scala 19:19]
  wire  top_reset; // @[SimTop.scala 19:19]
  wire  top_io_out_aw_ready; // @[SimTop.scala 19:19]
  wire  top_io_out_aw_valid; // @[SimTop.scala 19:19]
  wire [31:0] top_io_out_aw_bits_addr; // @[SimTop.scala 19:19]
  wire  top_io_out_w_ready; // @[SimTop.scala 19:19]
  wire  top_io_out_w_valid; // @[SimTop.scala 19:19]
  wire [63:0] top_io_out_w_bits_data; // @[SimTop.scala 19:19]
  wire [7:0] top_io_out_w_bits_strb; // @[SimTop.scala 19:19]
  wire  top_io_out_w_bits_last; // @[SimTop.scala 19:19]
  wire  top_io_out_b_ready; // @[SimTop.scala 19:19]
  wire  top_io_out_b_valid; // @[SimTop.scala 19:19]
  wire  top_io_out_ar_ready; // @[SimTop.scala 19:19]
  wire  top_io_out_ar_valid; // @[SimTop.scala 19:19]
  wire [31:0] top_io_out_ar_bits_addr; // @[SimTop.scala 19:19]
  wire  top_io_out_r_ready; // @[SimTop.scala 19:19]
  wire  top_io_out_r_valid; // @[SimTop.scala 19:19]
  wire [63:0] top_io_out_r_bits_data; // @[SimTop.scala 19:19]
  wire  top_io_out_r_bits_last; // @[SimTop.scala 19:19]
  wire  top_io_imem_inst_valid; // @[SimTop.scala 19:19]
  wire  top_io_imem_inst_ready; // @[SimTop.scala 19:19]
  wire [31:0] top_io_imem_inst_addr; // @[SimTop.scala 19:19]
  wire [127:0] top_io_imem_inst_read; // @[SimTop.scala 19:19]
  wire  top_io_dmem_data_valid; // @[SimTop.scala 19:19]
  wire  top_io_dmem_data_ready; // @[SimTop.scala 19:19]
  wire  top_io_dmem_data_req; // @[SimTop.scala 19:19]
  wire [31:0] top_io_dmem_data_addr; // @[SimTop.scala 19:19]
  wire [7:0] top_io_dmem_data_strb; // @[SimTop.scala 19:19]
  wire [127:0] top_io_dmem_data_read; // @[SimTop.scala 19:19]
  wire [127:0] top_io_dmem_data_write; // @[SimTop.scala 19:19]
  Core core ( // @[SimTop.scala 15:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_inst_valid(core_io_imem_inst_valid),
    .io_imem_inst_ready(core_io_imem_inst_ready),
    .io_imem_inst_addr(core_io_imem_inst_addr),
    .io_imem_inst_read(core_io_imem_inst_read),
    .io_dmem_data_valid(core_io_dmem_data_valid),
    .io_dmem_data_ready(core_io_dmem_data_ready),
    .io_dmem_data_req(core_io_dmem_data_req),
    .io_dmem_data_addr(core_io_dmem_data_addr),
    .io_dmem_data_size(core_io_dmem_data_size),
    .io_dmem_data_strb(core_io_dmem_data_strb),
    .io_dmem_data_read(core_io_dmem_data_read),
    .io_dmem_data_write(core_io_dmem_data_write)
  );
  Icache icache ( // @[SimTop.scala 16:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_imem_inst_valid(icache_io_imem_inst_valid),
    .io_imem_inst_ready(icache_io_imem_inst_ready),
    .io_imem_inst_addr(icache_io_imem_inst_addr),
    .io_imem_inst_read(icache_io_imem_inst_read),
    .io_out_inst_valid(icache_io_out_inst_valid),
    .io_out_inst_ready(icache_io_out_inst_ready),
    .io_out_inst_addr(icache_io_out_inst_addr),
    .io_out_inst_read(icache_io_out_inst_read)
  );
  Dcache dcache ( // @[SimTop.scala 17:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_dmem_data_valid(dcache_io_dmem_data_valid),
    .io_dmem_data_ready(dcache_io_dmem_data_ready),
    .io_dmem_data_req(dcache_io_dmem_data_req),
    .io_dmem_data_addr(dcache_io_dmem_data_addr),
    .io_dmem_data_size(dcache_io_dmem_data_size),
    .io_dmem_data_strb(dcache_io_dmem_data_strb),
    .io_dmem_data_read(dcache_io_dmem_data_read),
    .io_dmem_data_write(dcache_io_dmem_data_write),
    .io_out_data_valid(dcache_io_out_data_valid),
    .io_out_data_ready(dcache_io_out_data_ready),
    .io_out_data_req(dcache_io_out_data_req),
    .io_out_data_addr(dcache_io_out_data_addr),
    .io_out_data_strb(dcache_io_out_data_strb),
    .io_out_data_read(dcache_io_out_data_read),
    .io_out_data_write(dcache_io_out_data_write)
  );
  AxiLite2Axi top ( // @[SimTop.scala 19:19]
    .clock(top_clock),
    .reset(top_reset),
    .io_out_aw_ready(top_io_out_aw_ready),
    .io_out_aw_valid(top_io_out_aw_valid),
    .io_out_aw_bits_addr(top_io_out_aw_bits_addr),
    .io_out_w_ready(top_io_out_w_ready),
    .io_out_w_valid(top_io_out_w_valid),
    .io_out_w_bits_data(top_io_out_w_bits_data),
    .io_out_w_bits_strb(top_io_out_w_bits_strb),
    .io_out_w_bits_last(top_io_out_w_bits_last),
    .io_out_b_ready(top_io_out_b_ready),
    .io_out_b_valid(top_io_out_b_valid),
    .io_out_ar_ready(top_io_out_ar_ready),
    .io_out_ar_valid(top_io_out_ar_valid),
    .io_out_ar_bits_addr(top_io_out_ar_bits_addr),
    .io_out_r_ready(top_io_out_r_ready),
    .io_out_r_valid(top_io_out_r_valid),
    .io_out_r_bits_data(top_io_out_r_bits_data),
    .io_out_r_bits_last(top_io_out_r_bits_last),
    .io_imem_inst_valid(top_io_imem_inst_valid),
    .io_imem_inst_ready(top_io_imem_inst_ready),
    .io_imem_inst_addr(top_io_imem_inst_addr),
    .io_imem_inst_read(top_io_imem_inst_read),
    .io_dmem_data_valid(top_io_dmem_data_valid),
    .io_dmem_data_ready(top_io_dmem_data_ready),
    .io_dmem_data_req(top_io_dmem_data_req),
    .io_dmem_data_addr(top_io_dmem_data_addr),
    .io_dmem_data_strb(top_io_dmem_data_strb),
    .io_dmem_data_read(top_io_dmem_data_read),
    .io_dmem_data_write(top_io_dmem_data_write)
  );
  assign io_uart_out_valid = 1'h0; // @[SimTop.scala 36:21]
  assign io_uart_out_ch = 8'h0; // @[SimTop.scala 37:18]
  assign io_uart_in_valid = 1'h0; // @[SimTop.scala 38:20]
  assign io_memAXI_0_aw_valid = top_io_out_aw_valid; // @[SimTop.scala 30:18]
  assign io_memAXI_0_aw_bits_addr = top_io_out_aw_bits_addr; // @[SimTop.scala 30:18]
  assign io_memAXI_0_aw_bits_prot = 3'h0; // @[SimTop.scala 30:18]
  assign io_memAXI_0_aw_bits_id = 4'h0; // @[SimTop.scala 30:18]
  assign io_memAXI_0_aw_bits_user = 1'h0; // @[SimTop.scala 30:18]
  assign io_memAXI_0_aw_bits_len = 8'h0; // @[SimTop.scala 30:18]
  assign io_memAXI_0_aw_bits_size = 3'h3; // @[SimTop.scala 30:18]
  assign io_memAXI_0_aw_bits_burst = 2'h1; // @[SimTop.scala 30:18]
  assign io_memAXI_0_aw_bits_lock = 1'h0; // @[SimTop.scala 30:18]
  assign io_memAXI_0_aw_bits_cache = 4'h2; // @[SimTop.scala 30:18]
  assign io_memAXI_0_aw_bits_qos = 4'h0; // @[SimTop.scala 30:18]
  assign io_memAXI_0_w_valid = top_io_out_w_valid; // @[SimTop.scala 31:18]
  assign io_memAXI_0_w_bits_data = top_io_out_w_bits_data; // @[SimTop.scala 31:18]
  assign io_memAXI_0_w_bits_strb = top_io_out_w_bits_strb; // @[SimTop.scala 31:18]
  assign io_memAXI_0_w_bits_last = 1'h1; // @[SimTop.scala 31:18]
  assign io_memAXI_0_b_ready = 1'h1; // @[SimTop.scala 32:18]
  assign io_memAXI_0_ar_valid = top_io_out_ar_valid; // @[SimTop.scala 33:18]
  assign io_memAXI_0_ar_bits_addr = top_io_out_ar_bits_addr; // @[SimTop.scala 33:18]
  assign io_memAXI_0_ar_bits_prot = 3'h0; // @[SimTop.scala 33:18]
  assign io_memAXI_0_ar_bits_id = 4'h0; // @[SimTop.scala 33:18]
  assign io_memAXI_0_ar_bits_user = 1'h0; // @[SimTop.scala 33:18]
  assign io_memAXI_0_ar_bits_len = 8'h1; // @[SimTop.scala 33:18]
  assign io_memAXI_0_ar_bits_size = 3'h3; // @[SimTop.scala 33:18]
  assign io_memAXI_0_ar_bits_burst = 2'h1; // @[SimTop.scala 33:18]
  assign io_memAXI_0_ar_bits_lock = 1'h0; // @[SimTop.scala 33:18]
  assign io_memAXI_0_ar_bits_cache = 4'h2; // @[SimTop.scala 33:18]
  assign io_memAXI_0_ar_bits_qos = 4'h0; // @[SimTop.scala 33:18]
  assign io_memAXI_0_r_ready = 1'h1; // @[SimTop.scala 34:18]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_imem_inst_ready = icache_io_imem_inst_ready; // @[SimTop.scala 21:17]
  assign core_io_imem_inst_read = icache_io_imem_inst_read; // @[SimTop.scala 21:17]
  assign core_io_dmem_data_ready = dcache_io_dmem_data_ready; // @[SimTop.scala 23:17]
  assign core_io_dmem_data_read = dcache_io_dmem_data_read; // @[SimTop.scala 23:17]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_imem_inst_valid = core_io_imem_inst_valid; // @[SimTop.scala 21:17]
  assign icache_io_imem_inst_addr = core_io_imem_inst_addr; // @[SimTop.scala 21:17]
  assign icache_io_out_inst_ready = top_io_imem_inst_ready; // @[SimTop.scala 22:17]
  assign icache_io_out_inst_read = top_io_imem_inst_read; // @[SimTop.scala 22:17]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_dmem_data_valid = core_io_dmem_data_valid; // @[SimTop.scala 23:17]
  assign dcache_io_dmem_data_req = core_io_dmem_data_req; // @[SimTop.scala 23:17]
  assign dcache_io_dmem_data_addr = core_io_dmem_data_addr; // @[SimTop.scala 23:17]
  assign dcache_io_dmem_data_size = core_io_dmem_data_size; // @[SimTop.scala 23:17]
  assign dcache_io_dmem_data_strb = core_io_dmem_data_strb; // @[SimTop.scala 23:17]
  assign dcache_io_dmem_data_write = core_io_dmem_data_write; // @[SimTop.scala 23:17]
  assign dcache_io_out_data_ready = top_io_dmem_data_ready; // @[SimTop.scala 24:17]
  assign dcache_io_out_data_read = top_io_dmem_data_read; // @[SimTop.scala 24:17]
  assign top_clock = clock;
  assign top_reset = reset;
  assign top_io_out_aw_ready = io_memAXI_0_aw_ready; // @[SimTop.scala 30:18]
  assign top_io_out_w_ready = io_memAXI_0_w_ready; // @[SimTop.scala 31:18]
  assign top_io_out_b_valid = io_memAXI_0_b_valid; // @[SimTop.scala 32:18]
  assign top_io_out_ar_ready = io_memAXI_0_ar_ready; // @[SimTop.scala 33:18]
  assign top_io_out_r_valid = io_memAXI_0_r_valid; // @[SimTop.scala 34:18]
  assign top_io_out_r_bits_data = io_memAXI_0_r_bits_data; // @[SimTop.scala 34:18]
  assign top_io_out_r_bits_last = io_memAXI_0_r_bits_last; // @[SimTop.scala 34:18]
  assign top_io_imem_inst_valid = icache_io_out_inst_valid; // @[SimTop.scala 22:17]
  assign top_io_imem_inst_addr = icache_io_out_inst_addr; // @[SimTop.scala 22:17]
  assign top_io_dmem_data_valid = dcache_io_out_data_valid; // @[SimTop.scala 24:17]
  assign top_io_dmem_data_req = dcache_io_out_data_req; // @[SimTop.scala 24:17]
  assign top_io_dmem_data_addr = dcache_io_out_data_addr; // @[SimTop.scala 24:17]
  assign top_io_dmem_data_strb = dcache_io_out_data_strb; // @[SimTop.scala 24:17]
  assign top_io_dmem_data_write = dcache_io_out_data_write; // @[SimTop.scala 24:17]
endmodule
